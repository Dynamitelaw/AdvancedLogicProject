
module pStore ( clk, clr, weightsIn, biasesIn, biasWriteEnable, sumOut );
  input [159:0] weightsIn;
  input [159:0] biasesIn;
  output [255:0] sumOut;
  input clk, clr, biasWriteEnable;
  wire   n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n322, n323, n324, n326, n327, n332, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n350, n351, n352,
         n354, n355, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n434, n442, n445, n447, n461, n462, n463, n464, n465, n466, n467,
         n468, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n551, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2299,
         n2300, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368;
  wire   [7:0] addWeight_0__add_s;
  wire   [7:0] addWeight_0__add_biasesStored;
  wire   [7:0] addWeight_1__add_s;
  wire   [7:0] addWeight_1__add_biasesStored;
  wire   [7:0] addWeight_2__add_s;
  wire   [7:0] addWeight_2__add_biasesStored;
  wire   [7:0] addWeight_3__add_s;
  wire   [7:0] addWeight_3__add_biasesStored;
  wire   [7:0] addWeight_4__add_s;
  wire   [7:0] addWeight_4__add_biasesStored;
  wire   [7:0] addWeight_5__add_s;
  wire   [7:0] addWeight_5__add_biasesStored;
  wire   [7:0] addWeight_6__add_s;
  wire   [7:0] addWeight_6__add_biasesStored;
  wire   [7:0] addWeight_7__add_s;
  wire   [7:0] addWeight_7__add_biasesStored;
  wire   [7:0] addWeight_8__add_s;
  wire   [7:0] addWeight_8__add_biasesStored;
  wire   [7:0] addWeight_9__add_s;
  wire   [7:0] addWeight_9__add_biasesStored;
  wire   [7:0] addWeight_10__add_s;
  wire   [7:0] addWeight_10__add_biasesStored;
  wire   [7:0] addWeight_11__add_s;
  wire   [7:0] addWeight_11__add_biasesStored;
  wire   [7:0] addWeight_12__add_s;
  wire   [7:0] addWeight_12__add_biasesStored;
  wire   [7:0] addWeight_13__add_s;
  wire   [7:0] addWeight_13__add_biasesStored;
  wire   [7:0] addWeight_14__add_s;
  wire   [7:0] addWeight_14__add_biasesStored;
  wire   [7:0] addWeight_15__add_s;
  wire   [7:0] addWeight_15__add_biasesStored;
  wire   [7:0] addWeight_16__add_s;
  wire   [7:0] addWeight_16__add_biasesStored;
  wire   [7:0] addWeight_17__add_s;
  wire   [7:0] addWeight_17__add_biasesStored;
  wire   [7:0] addWeight_18__add_s;
  wire   [7:0] addWeight_18__add_biasesStored;
  wire   [7:0] addWeight_19__add_s;
  wire   [7:0] addWeight_19__add_biasesStored;
  wire   [7:0] addWeight_20__add_s;
  wire   [7:0] addWeight_20__add_biasesStored;
  wire   [7:0] addWeight_21__add_s;
  wire   [7:0] addWeight_21__add_biasesStored;
  wire   [7:0] addWeight_22__add_s;
  wire   [7:0] addWeight_22__add_biasesStored;
  wire   [7:0] addWeight_23__add_s;
  wire   [7:0] addWeight_23__add_biasesStored;
  wire   [7:0] addWeight_24__add_s;
  wire   [7:0] addWeight_24__add_biasesStored;
  wire   [7:0] addWeight_25__add_s;
  wire   [7:0] addWeight_25__add_biasesStored;
  wire   [7:0] addWeight_26__add_s;
  wire   [7:0] addWeight_26__add_biasesStored;
  wire   [7:0] addWeight_27__add_s;
  wire   [7:0] addWeight_27__add_biasesStored;
  wire   [7:0] addWeight_28__add_s;
  wire   [7:0] addWeight_28__add_biasesStored;
  wire   [7:0] addWeight_29__add_s;
  wire   [7:0] addWeight_29__add_biasesStored;
  wire   [7:0] addWeight_30__add_s;
  wire   [7:0] addWeight_30__add_biasesStored;
  wire   [7:0] addWeight_31__add_s;
  wire   [7:0] addWeight_31__add_biasesStored;

  TLATXLTS addWeight_0__add_biasesStored_reg_0_ ( .G(n2368), .D(biasesIn[0]), 
        .Q(addWeight_0__add_biasesStored[0]) );
  TLATXLTS addWeight_0__add_biasesStored_reg_1_ ( .G(n2368), .D(biasesIn[1]), 
        .Q(addWeight_0__add_biasesStored[1]) );
  TLATXLTS addWeight_0__add_biasesStored_reg_2_ ( .G(n2368), .D(biasesIn[2]), 
        .Q(addWeight_0__add_biasesStored[2]) );
  TLATXLTS addWeight_0__add_biasesStored_reg_3_ ( .G(n2368), .D(biasesIn[3]), 
        .Q(addWeight_0__add_biasesStored[3]) );
  TLATXLTS addWeight_0__add_biasesStored_reg_7_ ( .G(n2300), .D(biasesIn[4]), 
        .Q(addWeight_0__add_biasesStored[7]) );
  TLATXLTS addWeight_1__add_biasesStored_reg_0_ ( .G(n2299), .D(biasesIn[5]), 
        .Q(addWeight_1__add_biasesStored[0]) );
  TLATXLTS addWeight_1__add_biasesStored_reg_1_ ( .G(n2300), .D(biasesIn[6]), 
        .Q(addWeight_1__add_biasesStored[1]) );
  TLATXLTS addWeight_1__add_biasesStored_reg_2_ ( .G(n2299), .D(biasesIn[7]), 
        .Q(addWeight_1__add_biasesStored[2]) );
  TLATXLTS addWeight_1__add_biasesStored_reg_3_ ( .G(n2367), .D(biasesIn[8]), 
        .Q(addWeight_1__add_biasesStored[3]) );
  TLATXLTS addWeight_1__add_biasesStored_reg_7_ ( .G(n2367), .D(biasesIn[9]), 
        .Q(addWeight_1__add_biasesStored[7]) );
  TLATXLTS addWeight_2__add_biasesStored_reg_0_ ( .G(n2367), .D(biasesIn[10]), 
        .Q(addWeight_2__add_biasesStored[0]) );
  TLATXLTS addWeight_2__add_biasesStored_reg_1_ ( .G(n2367), .D(biasesIn[11]), 
        .Q(addWeight_2__add_biasesStored[1]) );
  TLATXLTS addWeight_2__add_biasesStored_reg_2_ ( .G(n2366), .D(biasesIn[12]), 
        .Q(addWeight_2__add_biasesStored[2]) );
  TLATXLTS addWeight_2__add_biasesStored_reg_3_ ( .G(n2366), .D(biasesIn[13]), 
        .Q(addWeight_2__add_biasesStored[3]) );
  TLATXLTS addWeight_2__add_biasesStored_reg_7_ ( .G(n2366), .D(biasesIn[14]), 
        .Q(addWeight_2__add_biasesStored[7]) );
  TLATXLTS addWeight_3__add_biasesStored_reg_0_ ( .G(n2366), .D(biasesIn[15]), 
        .Q(addWeight_3__add_biasesStored[0]) );
  TLATXLTS addWeight_3__add_biasesStored_reg_1_ ( .G(n2365), .D(biasesIn[16]), 
        .Q(addWeight_3__add_biasesStored[1]) );
  TLATXLTS addWeight_3__add_biasesStored_reg_2_ ( .G(n2365), .D(biasesIn[17]), 
        .Q(addWeight_3__add_biasesStored[2]) );
  TLATXLTS addWeight_3__add_biasesStored_reg_3_ ( .G(n2365), .D(biasesIn[18]), 
        .Q(addWeight_3__add_biasesStored[3]) );
  TLATXLTS addWeight_3__add_biasesStored_reg_7_ ( .G(n2365), .D(biasesIn[19]), 
        .Q(addWeight_3__add_biasesStored[7]) );
  TLATXLTS addWeight_4__add_biasesStored_reg_0_ ( .G(n2364), .D(biasesIn[20]), 
        .Q(addWeight_4__add_biasesStored[0]) );
  TLATXLTS addWeight_4__add_biasesStored_reg_1_ ( .G(n2364), .D(biasesIn[21]), 
        .Q(addWeight_4__add_biasesStored[1]) );
  TLATXLTS addWeight_4__add_biasesStored_reg_2_ ( .G(n2364), .D(biasesIn[22]), 
        .Q(addWeight_4__add_biasesStored[2]) );
  TLATXLTS addWeight_4__add_biasesStored_reg_3_ ( .G(n2364), .D(biasesIn[23]), 
        .Q(addWeight_4__add_biasesStored[3]) );
  TLATXLTS addWeight_4__add_biasesStored_reg_7_ ( .G(n2363), .D(biasesIn[24]), 
        .Q(addWeight_4__add_biasesStored[7]) );
  TLATXLTS addWeight_5__add_biasesStored_reg_0_ ( .G(n2363), .D(biasesIn[25]), 
        .Q(addWeight_5__add_biasesStored[0]) );
  TLATXLTS addWeight_5__add_biasesStored_reg_1_ ( .G(n2363), .D(biasesIn[26]), 
        .Q(addWeight_5__add_biasesStored[1]) );
  TLATXLTS addWeight_5__add_biasesStored_reg_2_ ( .G(n2363), .D(biasesIn[27]), 
        .Q(addWeight_5__add_biasesStored[2]) );
  TLATXLTS addWeight_5__add_biasesStored_reg_3_ ( .G(n2362), .D(biasesIn[28]), 
        .Q(addWeight_5__add_biasesStored[3]) );
  TLATXLTS addWeight_5__add_biasesStored_reg_7_ ( .G(n2362), .D(biasesIn[29]), 
        .Q(addWeight_5__add_biasesStored[7]) );
  TLATXLTS addWeight_6__add_biasesStored_reg_0_ ( .G(n2362), .D(biasesIn[30]), 
        .Q(addWeight_6__add_biasesStored[0]) );
  TLATXLTS addWeight_6__add_biasesStored_reg_1_ ( .G(n2362), .D(biasesIn[31]), 
        .Q(addWeight_6__add_biasesStored[1]) );
  TLATXLTS addWeight_6__add_biasesStored_reg_2_ ( .G(n2361), .D(biasesIn[32]), 
        .Q(addWeight_6__add_biasesStored[2]) );
  TLATXLTS addWeight_6__add_biasesStored_reg_3_ ( .G(n2361), .D(biasesIn[33]), 
        .Q(addWeight_6__add_biasesStored[3]) );
  TLATXLTS addWeight_6__add_biasesStored_reg_7_ ( .G(n2361), .D(biasesIn[34]), 
        .Q(addWeight_6__add_biasesStored[7]) );
  TLATXLTS addWeight_7__add_biasesStored_reg_0_ ( .G(n2361), .D(biasesIn[35]), 
        .Q(addWeight_7__add_biasesStored[0]) );
  TLATXLTS addWeight_7__add_biasesStored_reg_1_ ( .G(n2360), .D(biasesIn[36]), 
        .Q(addWeight_7__add_biasesStored[1]) );
  TLATXLTS addWeight_7__add_biasesStored_reg_2_ ( .G(n2360), .D(biasesIn[37]), 
        .Q(addWeight_7__add_biasesStored[2]) );
  TLATXLTS addWeight_7__add_biasesStored_reg_3_ ( .G(n2360), .D(biasesIn[38]), 
        .Q(addWeight_7__add_biasesStored[3]) );
  TLATXLTS addWeight_7__add_biasesStored_reg_7_ ( .G(n2360), .D(biasesIn[39]), 
        .Q(addWeight_7__add_biasesStored[7]) );
  TLATXLTS addWeight_8__add_biasesStored_reg_0_ ( .G(n2359), .D(biasesIn[40]), 
        .Q(addWeight_8__add_biasesStored[0]) );
  TLATXLTS addWeight_8__add_biasesStored_reg_1_ ( .G(n2359), .D(biasesIn[41]), 
        .Q(addWeight_8__add_biasesStored[1]) );
  TLATXLTS addWeight_8__add_biasesStored_reg_2_ ( .G(n2359), .D(biasesIn[42]), 
        .Q(addWeight_8__add_biasesStored[2]) );
  TLATXLTS addWeight_8__add_biasesStored_reg_3_ ( .G(n2359), .D(biasesIn[43]), 
        .Q(addWeight_8__add_biasesStored[3]) );
  TLATXLTS addWeight_8__add_biasesStored_reg_7_ ( .G(n2358), .D(biasesIn[44]), 
        .Q(addWeight_8__add_biasesStored[7]) );
  TLATXLTS addWeight_9__add_biasesStored_reg_0_ ( .G(n2358), .D(biasesIn[45]), 
        .Q(addWeight_9__add_biasesStored[0]) );
  TLATXLTS addWeight_9__add_biasesStored_reg_1_ ( .G(n2358), .D(biasesIn[46]), 
        .Q(addWeight_9__add_biasesStored[1]) );
  TLATXLTS addWeight_9__add_biasesStored_reg_2_ ( .G(n2358), .D(biasesIn[47]), 
        .Q(addWeight_9__add_biasesStored[2]) );
  TLATXLTS addWeight_9__add_biasesStored_reg_3_ ( .G(n2357), .D(biasesIn[48]), 
        .Q(addWeight_9__add_biasesStored[3]) );
  TLATXLTS addWeight_9__add_biasesStored_reg_7_ ( .G(n2357), .D(biasesIn[49]), 
        .Q(addWeight_9__add_biasesStored[7]) );
  TLATXLTS addWeight_10__add_biasesStored_reg_0_ ( .G(n2357), .D(biasesIn[50]), 
        .Q(addWeight_10__add_biasesStored[0]) );
  TLATXLTS addWeight_10__add_biasesStored_reg_1_ ( .G(n2357), .D(biasesIn[51]), 
        .Q(addWeight_10__add_biasesStored[1]) );
  TLATXLTS addWeight_10__add_biasesStored_reg_2_ ( .G(n2356), .D(biasesIn[52]), 
        .Q(addWeight_10__add_biasesStored[2]) );
  TLATXLTS addWeight_10__add_biasesStored_reg_3_ ( .G(n2356), .D(biasesIn[53]), 
        .Q(addWeight_10__add_biasesStored[3]) );
  TLATXLTS addWeight_10__add_biasesStored_reg_7_ ( .G(n2356), .D(biasesIn[54]), 
        .Q(addWeight_10__add_biasesStored[7]) );
  TLATXLTS addWeight_11__add_biasesStored_reg_0_ ( .G(n2356), .D(biasesIn[55]), 
        .Q(addWeight_11__add_biasesStored[0]) );
  TLATXLTS addWeight_11__add_biasesStored_reg_1_ ( .G(n2355), .D(biasesIn[56]), 
        .Q(addWeight_11__add_biasesStored[1]) );
  TLATXLTS addWeight_11__add_biasesStored_reg_2_ ( .G(n2355), .D(biasesIn[57]), 
        .Q(addWeight_11__add_biasesStored[2]) );
  TLATXLTS addWeight_11__add_biasesStored_reg_3_ ( .G(n2355), .D(biasesIn[58]), 
        .Q(addWeight_11__add_biasesStored[3]) );
  TLATXLTS addWeight_11__add_biasesStored_reg_7_ ( .G(n2355), .D(biasesIn[59]), 
        .Q(addWeight_11__add_biasesStored[7]) );
  TLATXLTS addWeight_12__add_biasesStored_reg_0_ ( .G(n2354), .D(biasesIn[60]), 
        .Q(addWeight_12__add_biasesStored[0]) );
  TLATXLTS addWeight_12__add_biasesStored_reg_1_ ( .G(n2354), .D(biasesIn[61]), 
        .Q(addWeight_12__add_biasesStored[1]) );
  TLATXLTS addWeight_12__add_biasesStored_reg_2_ ( .G(n2354), .D(biasesIn[62]), 
        .Q(addWeight_12__add_biasesStored[2]) );
  TLATXLTS addWeight_12__add_biasesStored_reg_3_ ( .G(n2354), .D(biasesIn[63]), 
        .Q(addWeight_12__add_biasesStored[3]) );
  TLATXLTS addWeight_12__add_biasesStored_reg_7_ ( .G(n2353), .D(biasesIn[64]), 
        .Q(addWeight_12__add_biasesStored[7]) );
  TLATXLTS addWeight_13__add_biasesStored_reg_0_ ( .G(n2353), .D(biasesIn[65]), 
        .Q(addWeight_13__add_biasesStored[0]) );
  TLATXLTS addWeight_13__add_biasesStored_reg_1_ ( .G(n2353), .D(biasesIn[66]), 
        .Q(addWeight_13__add_biasesStored[1]) );
  TLATXLTS addWeight_13__add_biasesStored_reg_2_ ( .G(n2353), .D(biasesIn[67]), 
        .Q(addWeight_13__add_biasesStored[2]) );
  TLATXLTS addWeight_13__add_biasesStored_reg_3_ ( .G(n2352), .D(biasesIn[68]), 
        .Q(addWeight_13__add_biasesStored[3]) );
  TLATXLTS addWeight_13__add_biasesStored_reg_7_ ( .G(n2352), .D(biasesIn[69]), 
        .Q(addWeight_13__add_biasesStored[7]) );
  TLATXLTS addWeight_14__add_biasesStored_reg_0_ ( .G(n2352), .D(biasesIn[70]), 
        .Q(addWeight_14__add_biasesStored[0]) );
  TLATXLTS addWeight_14__add_biasesStored_reg_1_ ( .G(n2352), .D(biasesIn[71]), 
        .Q(addWeight_14__add_biasesStored[1]) );
  TLATXLTS addWeight_14__add_biasesStored_reg_2_ ( .G(n2351), .D(biasesIn[72]), 
        .Q(addWeight_14__add_biasesStored[2]) );
  TLATXLTS addWeight_14__add_biasesStored_reg_3_ ( .G(n2351), .D(biasesIn[73]), 
        .Q(addWeight_14__add_biasesStored[3]) );
  TLATXLTS addWeight_14__add_biasesStored_reg_7_ ( .G(n2351), .D(biasesIn[74]), 
        .Q(addWeight_14__add_biasesStored[7]) );
  TLATXLTS addWeight_15__add_biasesStored_reg_0_ ( .G(n2351), .D(biasesIn[75]), 
        .Q(addWeight_15__add_biasesStored[0]) );
  TLATXLTS addWeight_15__add_biasesStored_reg_1_ ( .G(n2350), .D(biasesIn[76]), 
        .Q(addWeight_15__add_biasesStored[1]) );
  TLATXLTS addWeight_15__add_biasesStored_reg_2_ ( .G(n2350), .D(biasesIn[77]), 
        .Q(addWeight_15__add_biasesStored[2]) );
  TLATXLTS addWeight_15__add_biasesStored_reg_3_ ( .G(n2350), .D(biasesIn[78]), 
        .Q(addWeight_15__add_biasesStored[3]) );
  TLATXLTS addWeight_15__add_biasesStored_reg_7_ ( .G(n2350), .D(biasesIn[79]), 
        .Q(addWeight_15__add_biasesStored[7]) );
  TLATXLTS addWeight_16__add_biasesStored_reg_0_ ( .G(n2349), .D(biasesIn[80]), 
        .Q(addWeight_16__add_biasesStored[0]) );
  TLATXLTS addWeight_16__add_biasesStored_reg_1_ ( .G(n2349), .D(biasesIn[81]), 
        .Q(addWeight_16__add_biasesStored[1]) );
  TLATXLTS addWeight_16__add_biasesStored_reg_2_ ( .G(n2349), .D(biasesIn[82]), 
        .Q(addWeight_16__add_biasesStored[2]) );
  TLATXLTS addWeight_16__add_biasesStored_reg_3_ ( .G(n2349), .D(biasesIn[83]), 
        .Q(addWeight_16__add_biasesStored[3]) );
  TLATXLTS addWeight_16__add_biasesStored_reg_7_ ( .G(n2348), .D(biasesIn[84]), 
        .Q(addWeight_16__add_biasesStored[7]) );
  TLATXLTS addWeight_17__add_biasesStored_reg_0_ ( .G(n2348), .D(biasesIn[85]), 
        .Q(addWeight_17__add_biasesStored[0]) );
  TLATXLTS addWeight_17__add_biasesStored_reg_1_ ( .G(n2348), .D(biasesIn[86]), 
        .Q(addWeight_17__add_biasesStored[1]) );
  TLATXLTS addWeight_17__add_biasesStored_reg_2_ ( .G(n2348), .D(biasesIn[87]), 
        .Q(addWeight_17__add_biasesStored[2]) );
  TLATXLTS addWeight_17__add_biasesStored_reg_3_ ( .G(n2347), .D(biasesIn[88]), 
        .Q(addWeight_17__add_biasesStored[3]) );
  TLATXLTS addWeight_17__add_biasesStored_reg_7_ ( .G(n2347), .D(biasesIn[89]), 
        .Q(addWeight_17__add_biasesStored[7]) );
  TLATXLTS addWeight_18__add_biasesStored_reg_0_ ( .G(n2347), .D(biasesIn[90]), 
        .Q(addWeight_18__add_biasesStored[0]) );
  TLATXLTS addWeight_18__add_biasesStored_reg_1_ ( .G(n2347), .D(biasesIn[91]), 
        .Q(addWeight_18__add_biasesStored[1]) );
  TLATXLTS addWeight_18__add_biasesStored_reg_2_ ( .G(n2346), .D(biasesIn[92]), 
        .Q(addWeight_18__add_biasesStored[2]) );
  TLATXLTS addWeight_18__add_biasesStored_reg_3_ ( .G(n2346), .D(biasesIn[93]), 
        .Q(addWeight_18__add_biasesStored[3]) );
  TLATXLTS addWeight_18__add_biasesStored_reg_7_ ( .G(n2346), .D(biasesIn[94]), 
        .Q(addWeight_18__add_biasesStored[7]) );
  TLATXLTS addWeight_19__add_biasesStored_reg_0_ ( .G(n2346), .D(biasesIn[95]), 
        .Q(addWeight_19__add_biasesStored[0]) );
  TLATXLTS addWeight_19__add_biasesStored_reg_1_ ( .G(n2345), .D(biasesIn[96]), 
        .Q(addWeight_19__add_biasesStored[1]) );
  TLATXLTS addWeight_19__add_biasesStored_reg_2_ ( .G(n2345), .D(biasesIn[97]), 
        .Q(addWeight_19__add_biasesStored[2]) );
  TLATXLTS addWeight_19__add_biasesStored_reg_3_ ( .G(n2345), .D(biasesIn[98]), 
        .Q(addWeight_19__add_biasesStored[3]) );
  TLATXLTS addWeight_19__add_biasesStored_reg_7_ ( .G(n2345), .D(biasesIn[99]), 
        .Q(addWeight_19__add_biasesStored[7]) );
  TLATXLTS addWeight_20__add_biasesStored_reg_0_ ( .G(n2344), .D(biasesIn[100]), .Q(addWeight_20__add_biasesStored[0]) );
  TLATXLTS addWeight_20__add_biasesStored_reg_1_ ( .G(n2344), .D(biasesIn[101]), .Q(addWeight_20__add_biasesStored[1]) );
  TLATXLTS addWeight_20__add_biasesStored_reg_2_ ( .G(n2344), .D(biasesIn[102]), .Q(addWeight_20__add_biasesStored[2]) );
  TLATXLTS addWeight_20__add_biasesStored_reg_3_ ( .G(n2344), .D(biasesIn[103]), .Q(addWeight_20__add_biasesStored[3]) );
  TLATXLTS addWeight_20__add_biasesStored_reg_7_ ( .G(n2343), .D(biasesIn[104]), .Q(addWeight_20__add_biasesStored[7]) );
  TLATXLTS addWeight_21__add_biasesStored_reg_0_ ( .G(n2343), .D(biasesIn[105]), .Q(addWeight_21__add_biasesStored[0]) );
  TLATXLTS addWeight_21__add_biasesStored_reg_1_ ( .G(n2343), .D(biasesIn[106]), .Q(addWeight_21__add_biasesStored[1]) );
  TLATXLTS addWeight_21__add_biasesStored_reg_2_ ( .G(n2343), .D(biasesIn[107]), .Q(addWeight_21__add_biasesStored[2]) );
  TLATXLTS addWeight_21__add_biasesStored_reg_3_ ( .G(n2342), .D(biasesIn[108]), .Q(addWeight_21__add_biasesStored[3]) );
  TLATXLTS addWeight_21__add_biasesStored_reg_7_ ( .G(n2342), .D(biasesIn[109]), .Q(addWeight_21__add_biasesStored[7]) );
  TLATXLTS addWeight_22__add_biasesStored_reg_0_ ( .G(n2342), .D(biasesIn[110]), .Q(addWeight_22__add_biasesStored[0]) );
  TLATXLTS addWeight_22__add_biasesStored_reg_1_ ( .G(n2342), .D(biasesIn[111]), .Q(addWeight_22__add_biasesStored[1]) );
  TLATXLTS addWeight_22__add_biasesStored_reg_2_ ( .G(n2341), .D(biasesIn[112]), .Q(addWeight_22__add_biasesStored[2]) );
  TLATXLTS addWeight_22__add_biasesStored_reg_3_ ( .G(n2341), .D(biasesIn[113]), .Q(addWeight_22__add_biasesStored[3]) );
  TLATXLTS addWeight_22__add_biasesStored_reg_7_ ( .G(n2341), .D(biasesIn[114]), .Q(addWeight_22__add_biasesStored[7]) );
  TLATXLTS addWeight_23__add_biasesStored_reg_0_ ( .G(n2341), .D(biasesIn[115]), .Q(addWeight_23__add_biasesStored[0]) );
  TLATXLTS addWeight_23__add_biasesStored_reg_1_ ( .G(n2340), .D(biasesIn[116]), .Q(addWeight_23__add_biasesStored[1]) );
  TLATXLTS addWeight_23__add_biasesStored_reg_2_ ( .G(n2340), .D(biasesIn[117]), .Q(addWeight_23__add_biasesStored[2]) );
  TLATXLTS addWeight_23__add_biasesStored_reg_3_ ( .G(n2340), .D(biasesIn[118]), .Q(addWeight_23__add_biasesStored[3]) );
  TLATXLTS addWeight_23__add_biasesStored_reg_7_ ( .G(n2340), .D(biasesIn[119]), .Q(addWeight_23__add_biasesStored[7]) );
  TLATXLTS addWeight_24__add_biasesStored_reg_0_ ( .G(n2339), .D(biasesIn[120]), .Q(addWeight_24__add_biasesStored[0]) );
  TLATXLTS addWeight_24__add_biasesStored_reg_1_ ( .G(n2339), .D(biasesIn[121]), .Q(addWeight_24__add_biasesStored[1]) );
  TLATXLTS addWeight_24__add_biasesStored_reg_2_ ( .G(n2339), .D(biasesIn[122]), .Q(addWeight_24__add_biasesStored[2]) );
  TLATXLTS addWeight_24__add_biasesStored_reg_3_ ( .G(n2339), .D(biasesIn[123]), .Q(addWeight_24__add_biasesStored[3]) );
  TLATXLTS addWeight_24__add_biasesStored_reg_7_ ( .G(n2338), .D(biasesIn[124]), .Q(addWeight_24__add_biasesStored[7]) );
  TLATXLTS addWeight_25__add_biasesStored_reg_0_ ( .G(n2338), .D(biasesIn[125]), .Q(addWeight_25__add_biasesStored[0]) );
  TLATXLTS addWeight_25__add_biasesStored_reg_1_ ( .G(n2338), .D(biasesIn[126]), .Q(addWeight_25__add_biasesStored[1]) );
  TLATXLTS addWeight_25__add_biasesStored_reg_2_ ( .G(n2338), .D(biasesIn[127]), .Q(addWeight_25__add_biasesStored[2]) );
  TLATXLTS addWeight_25__add_biasesStored_reg_3_ ( .G(n2337), .D(biasesIn[128]), .Q(addWeight_25__add_biasesStored[3]) );
  TLATXLTS addWeight_25__add_biasesStored_reg_7_ ( .G(n2337), .D(biasesIn[129]), .Q(addWeight_25__add_biasesStored[7]) );
  TLATXLTS addWeight_26__add_biasesStored_reg_0_ ( .G(n2337), .D(biasesIn[130]), .Q(addWeight_26__add_biasesStored[0]) );
  TLATXLTS addWeight_26__add_biasesStored_reg_1_ ( .G(n2337), .D(biasesIn[131]), .Q(addWeight_26__add_biasesStored[1]) );
  TLATXLTS addWeight_26__add_biasesStored_reg_2_ ( .G(n2336), .D(biasesIn[132]), .Q(addWeight_26__add_biasesStored[2]) );
  TLATXLTS addWeight_26__add_biasesStored_reg_3_ ( .G(n2336), .D(biasesIn[133]), .Q(addWeight_26__add_biasesStored[3]) );
  TLATXLTS addWeight_26__add_biasesStored_reg_7_ ( .G(n2336), .D(biasesIn[134]), .Q(addWeight_26__add_biasesStored[7]) );
  TLATXLTS addWeight_27__add_biasesStored_reg_0_ ( .G(n2336), .D(biasesIn[135]), .Q(addWeight_27__add_biasesStored[0]) );
  TLATXLTS addWeight_27__add_biasesStored_reg_1_ ( .G(n2335), .D(biasesIn[136]), .Q(addWeight_27__add_biasesStored[1]) );
  TLATXLTS addWeight_27__add_biasesStored_reg_2_ ( .G(n2335), .D(biasesIn[137]), .Q(addWeight_27__add_biasesStored[2]) );
  TLATXLTS addWeight_27__add_biasesStored_reg_3_ ( .G(n2335), .D(biasesIn[138]), .Q(addWeight_27__add_biasesStored[3]) );
  TLATXLTS addWeight_27__add_biasesStored_reg_7_ ( .G(n2335), .D(biasesIn[139]), .Q(addWeight_27__add_biasesStored[7]) );
  TLATXLTS addWeight_28__add_biasesStored_reg_0_ ( .G(n2334), .D(biasesIn[140]), .Q(addWeight_28__add_biasesStored[0]) );
  TLATXLTS addWeight_28__add_biasesStored_reg_1_ ( .G(n2334), .D(biasesIn[141]), .Q(addWeight_28__add_biasesStored[1]) );
  TLATXLTS addWeight_28__add_biasesStored_reg_2_ ( .G(n2334), .D(biasesIn[142]), .Q(addWeight_28__add_biasesStored[2]) );
  TLATXLTS addWeight_28__add_biasesStored_reg_3_ ( .G(n2334), .D(biasesIn[143]), .Q(addWeight_28__add_biasesStored[3]) );
  TLATXLTS addWeight_28__add_biasesStored_reg_7_ ( .G(n2333), .D(biasesIn[144]), .Q(addWeight_28__add_biasesStored[7]) );
  TLATXLTS addWeight_29__add_biasesStored_reg_0_ ( .G(n2333), .D(biasesIn[145]), .Q(addWeight_29__add_biasesStored[0]) );
  TLATXLTS addWeight_29__add_biasesStored_reg_1_ ( .G(n2333), .D(biasesIn[146]), .Q(addWeight_29__add_biasesStored[1]) );
  TLATXLTS addWeight_29__add_biasesStored_reg_2_ ( .G(n2333), .D(biasesIn[147]), .Q(addWeight_29__add_biasesStored[2]) );
  TLATXLTS addWeight_29__add_biasesStored_reg_3_ ( .G(n2136), .D(biasesIn[148]), .Q(addWeight_29__add_biasesStored[3]) );
  TLATXLTS addWeight_29__add_biasesStored_reg_7_ ( .G(n2076), .D(biasesIn[149]), .Q(addWeight_29__add_biasesStored[7]) );
  TLATXLTS addWeight_30__add_biasesStored_reg_0_ ( .G(biasWriteEnable), .D(
        biasesIn[150]), .Q(addWeight_30__add_biasesStored[0]) );
  TLATXLTS addWeight_30__add_biasesStored_reg_1_ ( .G(biasWriteEnable), .D(
        biasesIn[151]), .Q(addWeight_30__add_biasesStored[1]) );
  TLATXLTS addWeight_30__add_biasesStored_reg_2_ ( .G(n2332), .D(biasesIn[152]), .Q(addWeight_30__add_biasesStored[2]) );
  TLATXLTS addWeight_30__add_biasesStored_reg_3_ ( .G(n2332), .D(biasesIn[153]), .Q(addWeight_30__add_biasesStored[3]) );
  TLATXLTS addWeight_30__add_biasesStored_reg_7_ ( .G(n2332), .D(biasesIn[154]), .Q(addWeight_30__add_biasesStored[7]) );
  TLATXLTS addWeight_31__add_biasesStored_reg_0_ ( .G(n2332), .D(biasesIn[155]), .Q(addWeight_31__add_biasesStored[0]) );
  TLATXLTS addWeight_31__add_biasesStored_reg_1_ ( .G(n2331), .D(biasesIn[156]), .Q(addWeight_31__add_biasesStored[1]) );
  TLATXLTS addWeight_31__add_biasesStored_reg_2_ ( .G(n2331), .D(biasesIn[157]), .Q(addWeight_31__add_biasesStored[2]) );
  TLATXLTS addWeight_31__add_biasesStored_reg_3_ ( .G(n2331), .D(biasesIn[158]), .Q(addWeight_31__add_biasesStored[3]) );
  TLATXLTS addWeight_31__add_biasesStored_reg_7_ ( .G(n2331), .D(biasesIn[159]), .Q(addWeight_31__add_biasesStored[7]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_6_ ( .D(addWeight_25__add_s[6]), .CK(clk), .SN(n257), .RN(n258), .Q(sumOut[206]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_5_ ( .D(addWeight_25__add_s[5]), .CK(clk), .SN(n257), .RN(n258), .Q(sumOut[205]) );
  DFFSRHQX4TS addWeight_3__add_S_reg_7_ ( .D(addWeight_3__add_s[7]), .CK(clk), 
        .SN(n37), .RN(n38), .Q(sumOut[31]) );
  DFFSRHQX4TS addWeight_4__add_S_reg_7_ ( .D(addWeight_4__add_s[7]), .CK(clk), 
        .SN(n47), .RN(n48), .Q(sumOut[39]) );
  DFFSRHQX4TS addWeight_5__add_S_reg_7_ ( .D(addWeight_5__add_s[7]), .CK(clk), 
        .SN(n57), .RN(n58), .Q(sumOut[47]) );
  DFFSRHQX4TS addWeight_6__add_S_reg_7_ ( .D(addWeight_6__add_s[7]), .CK(clk), 
        .SN(n67), .RN(n68), .Q(sumOut[55]) );
  DFFSRHQX4TS addWeight_7__add_S_reg_7_ ( .D(addWeight_7__add_s[7]), .CK(clk), 
        .SN(n77), .RN(n78), .Q(sumOut[63]) );
  DFFSRHQX4TS addWeight_8__add_S_reg_7_ ( .D(addWeight_8__add_s[7]), .CK(clk), 
        .SN(n87), .RN(n88), .Q(sumOut[71]) );
  DFFSRHQX4TS addWeight_9__add_S_reg_7_ ( .D(addWeight_9__add_s[7]), .CK(clk), 
        .SN(n97), .RN(n98), .Q(sumOut[79]) );
  DFFSRHQX4TS addWeight_13__add_S_reg_7_ ( .D(addWeight_13__add_s[7]), .CK(clk), .SN(n137), .RN(n138), .Q(sumOut[111]) );
  DFFSRHQX4TS addWeight_14__add_S_reg_7_ ( .D(addWeight_14__add_s[7]), .CK(clk), .SN(n147), .RN(n148), .Q(sumOut[119]) );
  DFFSRHQX4TS addWeight_15__add_S_reg_7_ ( .D(addWeight_15__add_s[7]), .CK(clk), .SN(n157), .RN(n158), .Q(sumOut[127]) );
  DFFSRHQX4TS addWeight_16__add_S_reg_7_ ( .D(addWeight_16__add_s[7]), .CK(clk), .SN(n167), .RN(n168), .Q(sumOut[135]) );
  DFFSRHQX4TS addWeight_17__add_S_reg_7_ ( .D(addWeight_17__add_s[7]), .CK(clk), .SN(n177), .RN(n178), .Q(sumOut[143]) );
  DFFSRHQX4TS addWeight_18__add_S_reg_7_ ( .D(addWeight_18__add_s[7]), .CK(clk), .SN(n187), .RN(n188), .Q(sumOut[151]) );
  DFFSRHQX4TS addWeight_19__add_S_reg_7_ ( .D(addWeight_19__add_s[7]), .CK(clk), .SN(n197), .RN(n198), .Q(sumOut[159]) );
  DFFSRHQX4TS addWeight_20__add_S_reg_7_ ( .D(addWeight_20__add_s[7]), .CK(clk), .SN(n207), .RN(n208), .Q(sumOut[167]) );
  DFFSRHQX4TS addWeight_21__add_S_reg_7_ ( .D(addWeight_21__add_s[7]), .CK(clk), .SN(n217), .RN(n218), .Q(sumOut[175]) );
  DFFSRHQX4TS addWeight_22__add_S_reg_7_ ( .D(addWeight_22__add_s[7]), .CK(clk), .SN(n227), .RN(n228), .Q(sumOut[183]) );
  DFFSRHQX4TS addWeight_23__add_S_reg_7_ ( .D(addWeight_23__add_s[7]), .CK(clk), .SN(n237), .RN(n238), .Q(sumOut[191]) );
  DFFSRHQX4TS addWeight_24__add_S_reg_7_ ( .D(addWeight_24__add_s[7]), .CK(clk), .SN(n247), .RN(n248), .Q(sumOut[199]) );
  DFFSRHQX4TS addWeight_30__add_S_reg_7_ ( .D(addWeight_30__add_s[7]), .CK(clk), .SN(n307), .RN(n308), .Q(sumOut[247]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_3_ ( .D(addWeight_25__add_s[3]), .CK(clk), .SN(n255), .RN(n256), .Q(sumOut[203]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_7_ ( .D(addWeight_11__add_s[7]), .CK(clk), .SN(n117), .RN(n118), .Q(sumOut[95]) );
  DFFSRHQX4TS addWeight_1__add_S_reg_7_ ( .D(addWeight_1__add_s[7]), .CK(clk), 
        .SN(n17), .RN(n18), .Q(sumOut[15]) );
  DFFSRHQX4TS addWeight_0__add_S_reg_7_ ( .D(addWeight_0__add_s[7]), .CK(clk), 
        .SN(n7), .RN(n8), .Q(sumOut[7]) );
  DFFSRHQX4TS addWeight_1__add_S_reg_6_ ( .D(addWeight_1__add_s[6]), .CK(clk), 
        .SN(n17), .RN(n18), .Q(sumOut[14]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_5_ ( .D(addWeight_2__add_s[5]), .CK(clk), 
        .SN(n27), .RN(n28), .Q(sumOut[21]) );
  DFFSRHQX4TS addWeight_20__add_S_reg_6_ ( .D(addWeight_20__add_s[6]), .CK(clk), .SN(n207), .RN(n208), .Q(sumOut[166]) );
  DFFSRHQX4TS addWeight_21__add_S_reg_6_ ( .D(addWeight_21__add_s[6]), .CK(clk), .SN(n217), .RN(n218), .Q(sumOut[174]) );
  DFFSRHQX4TS addWeight_22__add_S_reg_6_ ( .D(addWeight_22__add_s[6]), .CK(clk), .SN(n227), .RN(n228), .Q(sumOut[182]) );
  DFFSRHQX4TS addWeight_23__add_S_reg_6_ ( .D(addWeight_23__add_s[6]), .CK(clk), .SN(n237), .RN(n238), .Q(sumOut[190]) );
  DFFSRHQX4TS addWeight_24__add_S_reg_6_ ( .D(addWeight_24__add_s[6]), .CK(clk), .SN(n247), .RN(n248), .Q(sumOut[198]) );
  DFFSRHQX4TS addWeight_30__add_S_reg_6_ ( .D(addWeight_30__add_s[6]), .CK(clk), .SN(n307), .RN(n308), .Q(sumOut[246]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_2_ ( .D(addWeight_29__add_s[2]), .CK(clk), .SN(n293), .RN(n294), .Q(n2374) );
  DFFSRHQX4TS addWeight_0__add_S_reg_3_ ( .D(addWeight_0__add_s[3]), .CK(clk), 
        .SN(n5), .RN(n6), .Q(n2447) );
  DFFSRHQX4TS addWeight_31__add_S_reg_7_ ( .D(addWeight_31__add_s[7]), .CK(clk), .SN(n317), .RN(n318), .Q(sumOut[255]) );
  DFFSRHQX4TS addWeight_30__add_S_reg_5_ ( .D(addWeight_30__add_s[5]), .CK(clk), .SN(n307), .RN(n308), .Q(sumOut[245]) );
  DFFSRHQX4TS addWeight_24__add_S_reg_5_ ( .D(addWeight_24__add_s[5]), .CK(clk), .SN(n247), .RN(n248), .Q(sumOut[197]) );
  DFFSRHQX4TS addWeight_23__add_S_reg_5_ ( .D(addWeight_23__add_s[5]), .CK(clk), .SN(n237), .RN(n238), .Q(sumOut[189]) );
  DFFSRHQX4TS addWeight_22__add_S_reg_5_ ( .D(addWeight_22__add_s[5]), .CK(clk), .SN(n227), .RN(n228), .Q(sumOut[181]) );
  DFFSRHQX4TS addWeight_21__add_S_reg_5_ ( .D(addWeight_21__add_s[5]), .CK(clk), .SN(n217), .RN(n218), .Q(sumOut[173]) );
  DFFSRHQX4TS addWeight_20__add_S_reg_5_ ( .D(addWeight_20__add_s[5]), .CK(clk), .SN(n207), .RN(n208), .Q(sumOut[165]) );
  DFFSRHQX4TS addWeight_19__add_S_reg_5_ ( .D(addWeight_19__add_s[5]), .CK(clk), .SN(n197), .RN(n198), .Q(sumOut[157]) );
  DFFSRHQX4TS addWeight_19__add_S_reg_3_ ( .D(addWeight_19__add_s[3]), .CK(clk), .SN(n195), .RN(n196), .Q(n2395) );
  DFFSRHQX4TS addWeight_20__add_S_reg_3_ ( .D(addWeight_20__add_s[3]), .CK(clk), .SN(n205), .RN(n206), .Q(n2392) );
  DFFSRHQX4TS addWeight_21__add_S_reg_3_ ( .D(addWeight_21__add_s[3]), .CK(clk), .SN(n215), .RN(n216), .Q(n2390) );
  DFFSRHQX4TS addWeight_22__add_S_reg_3_ ( .D(addWeight_22__add_s[3]), .CK(clk), .SN(n225), .RN(n226), .Q(n2388) );
  DFFSRHQX4TS addWeight_23__add_S_reg_3_ ( .D(addWeight_23__add_s[3]), .CK(clk), .SN(n235), .RN(n236), .Q(n2386) );
  DFFSRHQX4TS addWeight_24__add_S_reg_3_ ( .D(addWeight_24__add_s[3]), .CK(clk), .SN(n245), .RN(n246), .Q(n2383) );
  DFFSRHQX4TS addWeight_30__add_S_reg_3_ ( .D(addWeight_30__add_s[3]), .CK(clk), .SN(n305), .RN(n306), .Q(n2371) );
  DFFSRHQX4TS addWeight_3__add_S_reg_3_ ( .D(addWeight_3__add_s[3]), .CK(clk), 
        .SN(n35), .RN(n36), .Q(n2440) );
  DFFSRHQX4TS addWeight_4__add_S_reg_3_ ( .D(addWeight_4__add_s[3]), .CK(clk), 
        .SN(n45), .RN(n46), .Q(n2437) );
  DFFSRHQX4TS addWeight_5__add_S_reg_3_ ( .D(addWeight_5__add_s[3]), .CK(clk), 
        .SN(n55), .RN(n56), .Q(n2434) );
  DFFSRHQX4TS addWeight_6__add_S_reg_3_ ( .D(addWeight_6__add_s[3]), .CK(clk), 
        .SN(n65), .RN(n66), .Q(n2431) );
  DFFSRHQX4TS addWeight_7__add_S_reg_3_ ( .D(addWeight_7__add_s[3]), .CK(clk), 
        .SN(n75), .RN(n76), .Q(n2428) );
  DFFSRHQX4TS addWeight_8__add_S_reg_3_ ( .D(addWeight_8__add_s[3]), .CK(clk), 
        .SN(n85), .RN(n86), .Q(n2425) );
  DFFSRHQX4TS addWeight_9__add_S_reg_3_ ( .D(addWeight_9__add_s[3]), .CK(clk), 
        .SN(n95), .RN(n96), .Q(n2422) );
  DFFSRHQX4TS addWeight_13__add_S_reg_3_ ( .D(addWeight_13__add_s[3]), .CK(clk), .SN(n135), .RN(n136), .Q(n2411) );
  DFFSRHQX4TS addWeight_14__add_S_reg_3_ ( .D(addWeight_14__add_s[3]), .CK(clk), .SN(n145), .RN(n146), .Q(n2408) );
  DFFSRHQX4TS addWeight_15__add_S_reg_3_ ( .D(addWeight_15__add_s[3]), .CK(clk), .SN(n155), .RN(n156), .Q(n2405) );
  DFFSRHQX4TS addWeight_16__add_S_reg_3_ ( .D(addWeight_16__add_s[3]), .CK(clk), .SN(n165), .RN(n166), .Q(n2403) );
  DFFSRHQX4TS addWeight_17__add_S_reg_3_ ( .D(addWeight_17__add_s[3]), .CK(clk), .SN(n175), .RN(n176), .Q(n2400) );
  DFFSRHQX4TS addWeight_18__add_S_reg_3_ ( .D(addWeight_18__add_s[3]), .CK(clk), .SN(n185), .RN(n186), .Q(n2397) );
  DFFSRHQX4TS addWeight_10__add_S_reg_3_ ( .D(addWeight_10__add_s[3]), .CK(clk), .SN(n105), .RN(n106), .Q(n2420) );
  DFFSRHQX4TS addWeight_31__add_S_reg_3_ ( .D(addWeight_31__add_s[3]), .CK(clk), .SN(n315), .RN(n316), .Q(n2369) );
  DFFSRHQX4TS addWeight_1__add_S_reg_3_ ( .D(addWeight_1__add_s[3]), .CK(clk), 
        .SN(n15), .RN(n16), .Q(n2444) );
  DFFSRHQX4TS addWeight_11__add_S_reg_3_ ( .D(addWeight_11__add_s[3]), .CK(clk), .SN(n115), .RN(n116), .Q(n2417) );
  DFFSRHQX4TS addWeight_28__add_S_reg_3_ ( .D(addWeight_28__add_s[3]), .CK(clk), .SN(n285), .RN(n286), .Q(n2377) );
  DFFSRHQX4TS addWeight_12__add_S_reg_3_ ( .D(addWeight_12__add_s[3]), .CK(clk), .SN(n125), .RN(n126), .Q(n2414) );
  DFFSRHQX4TS addWeight_1__add_S_reg_2_ ( .D(addWeight_1__add_s[2]), .CK(clk), 
        .SN(n13), .RN(n14), .Q(sumOut[10]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_2_ ( .D(addWeight_11__add_s[2]), .CK(clk), .SN(n113), .RN(n114), .Q(sumOut[90]) );
  DFFSRHQX4TS addWeight_28__add_S_reg_2_ ( .D(addWeight_28__add_s[2]), .CK(clk), .SN(n283), .RN(n284), .Q(sumOut[226]) );
  DFFSRHQX4TS addWeight_12__add_S_reg_2_ ( .D(addWeight_12__add_s[2]), .CK(clk), .SN(n123), .RN(n124), .Q(sumOut[98]) );
  DFFSRHQX4TS addWeight_0__add_S_reg_2_ ( .D(addWeight_0__add_s[2]), .CK(clk), 
        .SN(n3), .RN(n4), .Q(sumOut[2]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_2_ ( .D(addWeight_2__add_s[2]), .CK(clk), 
        .SN(n23), .RN(n24), .Q(sumOut[18]) );
  DFFSRHQX4TS addWeight_10__add_S_reg_2_ ( .D(addWeight_10__add_s[2]), .CK(clk), .SN(n103), .RN(n104), .Q(n2421) );
  DFFSRHQX4TS addWeight_19__add_S_reg_2_ ( .D(addWeight_19__add_s[2]), .CK(clk), .SN(n193), .RN(n194), .Q(n2396) );
  DFFSRHQX4TS addWeight_20__add_S_reg_2_ ( .D(addWeight_20__add_s[2]), .CK(clk), .SN(n203), .RN(n204), .Q(sumOut[162]) );
  DFFSRHQX4TS addWeight_21__add_S_reg_2_ ( .D(addWeight_21__add_s[2]), .CK(clk), .SN(n213), .RN(n214), .Q(sumOut[170]) );
  DFFSRHQX4TS addWeight_22__add_S_reg_2_ ( .D(addWeight_22__add_s[2]), .CK(clk), .SN(n223), .RN(n224), .Q(sumOut[178]) );
  DFFSRHQX4TS addWeight_23__add_S_reg_2_ ( .D(addWeight_23__add_s[2]), .CK(clk), .SN(n233), .RN(n234), .Q(sumOut[186]) );
  DFFSRHQX4TS addWeight_24__add_S_reg_2_ ( .D(addWeight_24__add_s[2]), .CK(clk), .SN(n243), .RN(n244), .Q(sumOut[194]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_2_ ( .D(addWeight_25__add_s[2]), .CK(clk), .SN(n253), .RN(n254), .Q(n2380) );
  DFFSRHQX4TS addWeight_27__add_S_reg_2_ ( .D(addWeight_27__add_s[2]), .CK(clk), .SN(n273), .RN(n274), .Q(sumOut[218]) );
  DFFSRHQX4TS addWeight_30__add_S_reg_2_ ( .D(addWeight_30__add_s[2]), .CK(clk), .SN(n303), .RN(n304), .Q(sumOut[242]) );
  DFFSRHQX4TS addWeight_31__add_S_reg_2_ ( .D(addWeight_31__add_s[2]), .CK(clk), .SN(n313), .RN(n314), .Q(sumOut[250]) );
  DFFSRHQX4TS addWeight_28__add_S_reg_1_ ( .D(addWeight_28__add_s[1]), .CK(clk), .SN(n281), .RN(n282), .Q(sumOut[225]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_1_ ( .D(addWeight_11__add_s[1]), .CK(clk), .SN(n111), .RN(n112), .Q(n2418) );
  DFFSRHQX4TS addWeight_1__add_S_reg_1_ ( .D(addWeight_1__add_s[1]), .CK(clk), 
        .SN(n11), .RN(n12), .Q(n2445) );
  DFFSRHQX4TS addWeight_12__add_S_reg_1_ ( .D(addWeight_12__add_s[1]), .CK(clk), .SN(n121), .RN(n122), .Q(n2415) );
  DFFSRHQX4TS addWeight_26__add_S_reg_1_ ( .D(addWeight_26__add_s[1]), .CK(clk), .SN(n261), .RN(n262), .Q(sumOut[209]) );
  DFFSRHQX4TS addWeight_27__add_S_reg_5_ ( .D(addWeight_27__add_s[5]), .CK(clk), .SN(n277), .RN(n278), .Q(sumOut[221]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_1_ ( .D(addWeight_25__add_s[1]), .CK(clk), .SN(n251), .RN(n252), .Q(n2381) );
  DFFSRHQX4TS addWeight_29__add_S_reg_3_ ( .D(addWeight_29__add_s[3]), .CK(clk), .SN(n295), .RN(n296), .Q(n2373) );
  DFFSRHQX4TS addWeight_17__add_S_reg_1_ ( .D(addWeight_17__add_s[1]), .CK(clk), .SN(n171), .RN(n172), .Q(n2401) );
  DFFSRHQX4TS addWeight_8__add_S_reg_1_ ( .D(addWeight_8__add_s[1]), .CK(clk), 
        .SN(n81), .RN(n82), .Q(n2426) );
  DFFSRHQX4TS addWeight_6__add_S_reg_1_ ( .D(addWeight_6__add_s[1]), .CK(clk), 
        .SN(n61), .RN(n62), .Q(n2432) );
  DFFSRHQX4TS addWeight_9__add_S_reg_1_ ( .D(addWeight_9__add_s[1]), .CK(clk), 
        .SN(n91), .RN(n92), .Q(n2423) );
  DFFSRHQX4TS addWeight_15__add_S_reg_1_ ( .D(addWeight_15__add_s[1]), .CK(clk), .SN(n151), .RN(n152), .Q(n2406) );
  DFFSRHQX4TS addWeight_7__add_S_reg_1_ ( .D(addWeight_7__add_s[1]), .CK(clk), 
        .SN(n71), .RN(n72), .Q(n2429) );
  DFFSRHQX4TS addWeight_13__add_S_reg_1_ ( .D(addWeight_13__add_s[1]), .CK(clk), .SN(n131), .RN(n132), .Q(n2412) );
  DFFSRHQX4TS addWeight_14__add_S_reg_1_ ( .D(addWeight_14__add_s[1]), .CK(clk), .SN(n141), .RN(n142), .Q(n2409) );
  DFFSRHQX4TS addWeight_18__add_S_reg_1_ ( .D(addWeight_18__add_s[1]), .CK(clk), .SN(n181), .RN(n182), .Q(n2398) );
  DFFSRHQX4TS addWeight_4__add_S_reg_1_ ( .D(addWeight_4__add_s[1]), .CK(clk), 
        .SN(n41), .RN(n42), .Q(n2438) );
  DFFSRHQX4TS addWeight_5__add_S_reg_1_ ( .D(addWeight_5__add_s[1]), .CK(clk), 
        .SN(n51), .RN(n52), .Q(n2435) );
  DFFSRHQX4TS addWeight_3__add_S_reg_1_ ( .D(addWeight_3__add_s[1]), .CK(clk), 
        .SN(n31), .RN(n32), .Q(n2441) );
  DFFSRHQX4TS addWeight_16__add_S_reg_1_ ( .D(addWeight_16__add_s[1]), .CK(clk), .SN(n161), .RN(n162), .Q(n2404) );
  DFFSRHQX4TS addWeight_19__add_S_reg_1_ ( .D(addWeight_19__add_s[1]), .CK(clk), .SN(n191), .RN(n192), .Q(sumOut[153]) );
  DFFSRHQX4TS addWeight_20__add_S_reg_1_ ( .D(addWeight_20__add_s[1]), .CK(clk), .SN(n201), .RN(n202), .Q(n2393) );
  DFFSRHQX4TS addWeight_30__add_S_reg_1_ ( .D(addWeight_30__add_s[1]), .CK(clk), .SN(n301), .RN(n302), .Q(n2372) );
  DFFSRHQX4TS addWeight_23__add_S_reg_1_ ( .D(addWeight_23__add_s[1]), .CK(clk), .SN(n231), .RN(n232), .Q(n2387) );
  DFFSRHQX4TS addWeight_24__add_S_reg_1_ ( .D(addWeight_24__add_s[1]), .CK(clk), .SN(n241), .RN(n242), .Q(n2384) );
  DFFSRHQX4TS addWeight_22__add_S_reg_1_ ( .D(addWeight_22__add_s[1]), .CK(clk), .SN(n221), .RN(n222), .Q(n2389) );
  DFFSRHQX4TS addWeight_21__add_S_reg_1_ ( .D(addWeight_21__add_s[1]), .CK(clk), .SN(n211), .RN(n212), .Q(n2391) );
  DFFSRHQX4TS addWeight_26__add_S_reg_0_ ( .D(addWeight_26__add_s[0]), .CK(clk), .SN(n269), .RN(n270), .Q(sumOut[208]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_0_ ( .D(addWeight_25__add_s[0]), .CK(clk), .SN(n259), .RN(n260), .Q(n2382) );
  DFFSRHQX4TS addWeight_27__add_S_reg_0_ ( .D(addWeight_27__add_s[0]), .CK(clk), .SN(n279), .RN(n280), .Q(sumOut[216]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_1_ ( .D(addWeight_29__add_s[1]), .CK(clk), .SN(n291), .RN(n292), .Q(n2375) );
  DFFSRHQX4TS addWeight_0__add_S_reg_0_ ( .D(addWeight_0__add_s[0]), .CK(clk), 
        .SN(n9), .RN(n10), .Q(sumOut[0]) );
  DFFSRHQX4TS addWeight_17__add_S_reg_2_ ( .D(addWeight_17__add_s[2]), .CK(clk), .SN(n173), .RN(n174), .Q(sumOut[138]) );
  DFFSRHQX4TS addWeight_8__add_S_reg_2_ ( .D(addWeight_8__add_s[2]), .CK(clk), 
        .SN(n83), .RN(n84), .Q(sumOut[66]) );
  DFFSRHQX4TS addWeight_6__add_S_reg_2_ ( .D(addWeight_6__add_s[2]), .CK(clk), 
        .SN(n63), .RN(n64), .Q(sumOut[50]) );
  DFFSRHQX4TS addWeight_9__add_S_reg_2_ ( .D(addWeight_9__add_s[2]), .CK(clk), 
        .SN(n93), .RN(n94), .Q(sumOut[74]) );
  DFFSRHQX4TS addWeight_15__add_S_reg_2_ ( .D(addWeight_15__add_s[2]), .CK(clk), .SN(n153), .RN(n154), .Q(sumOut[122]) );
  DFFSRHQX4TS addWeight_7__add_S_reg_2_ ( .D(addWeight_7__add_s[2]), .CK(clk), 
        .SN(n73), .RN(n74), .Q(sumOut[58]) );
  DFFSRHQX4TS addWeight_13__add_S_reg_2_ ( .D(addWeight_13__add_s[2]), .CK(clk), .SN(n133), .RN(n134), .Q(sumOut[106]) );
  DFFSRHQX4TS addWeight_14__add_S_reg_2_ ( .D(addWeight_14__add_s[2]), .CK(clk), .SN(n143), .RN(n144), .Q(sumOut[114]) );
  DFFSRHQX4TS addWeight_18__add_S_reg_2_ ( .D(addWeight_18__add_s[2]), .CK(clk), .SN(n183), .RN(n184), .Q(sumOut[146]) );
  DFFSRHQX4TS addWeight_4__add_S_reg_2_ ( .D(addWeight_4__add_s[2]), .CK(clk), 
        .SN(n43), .RN(n44), .Q(sumOut[34]) );
  DFFSRHQX4TS addWeight_5__add_S_reg_2_ ( .D(addWeight_5__add_s[2]), .CK(clk), 
        .SN(n53), .RN(n54), .Q(sumOut[42]) );
  DFFSRHQX4TS addWeight_3__add_S_reg_2_ ( .D(addWeight_3__add_s[2]), .CK(clk), 
        .SN(n33), .RN(n34), .Q(sumOut[26]) );
  DFFSRHQX4TS addWeight_16__add_S_reg_2_ ( .D(addWeight_16__add_s[2]), .CK(clk), .SN(n163), .RN(n164), .Q(sumOut[130]) );
  DFFSRHQX4TS addWeight_31__add_S_reg_1_ ( .D(addWeight_31__add_s[1]), .CK(clk), .SN(n311), .RN(n312), .Q(n2370) );
  DFFSRHQX4TS addWeight_10__add_S_reg_1_ ( .D(addWeight_10__add_s[1]), .CK(clk), .SN(n101), .RN(n102), .Q(sumOut[81]) );
  DFFSRHQX4TS addWeight_25__add_S_reg_4_ ( .D(addWeight_25__add_s[4]), .CK(clk), .SN(n257), .RN(n258), .Q(sumOut[204]) );
  DFFSRHQX4TS addWeight_0__add_S_reg_1_ ( .D(addWeight_0__add_s[1]), .CK(clk), 
        .SN(n1), .RN(n2), .Q(n2448) );
  DFFSRHQX4TS addWeight_27__add_S_reg_1_ ( .D(addWeight_27__add_s[1]), .CK(clk), .SN(n271), .RN(n272), .Q(sumOut[217]) );
  DFFSRHQX4TS addWeight_10__add_S_reg_0_ ( .D(addWeight_10__add_s[0]), .CK(clk), .SN(n109), .RN(n110), .Q(sumOut[80]) );
  DFFSRHQX4TS addWeight_31__add_S_reg_0_ ( .D(addWeight_31__add_s[0]), .CK(clk), .SN(n319), .RN(n320), .Q(sumOut[248]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_0_ ( .D(addWeight_29__add_s[0]), .CK(clk), .SN(n299), .RN(n300), .Q(n2376) );
  DFFSRHQX4TS addWeight_17__add_S_reg_0_ ( .D(addWeight_17__add_s[0]), .CK(clk), .SN(n179), .RN(n180), .Q(n2402) );
  DFFSRHQX4TS addWeight_8__add_S_reg_0_ ( .D(addWeight_8__add_s[0]), .CK(clk), 
        .SN(n89), .RN(n90), .Q(n2427) );
  DFFSRHQX4TS addWeight_6__add_S_reg_0_ ( .D(addWeight_6__add_s[0]), .CK(clk), 
        .SN(n69), .RN(n70), .Q(n2433) );
  DFFSRHQX4TS addWeight_9__add_S_reg_0_ ( .D(addWeight_9__add_s[0]), .CK(clk), 
        .SN(n99), .RN(n100), .Q(n2424) );
  DFFSRHQX4TS addWeight_15__add_S_reg_0_ ( .D(addWeight_15__add_s[0]), .CK(clk), .SN(n159), .RN(n160), .Q(n2407) );
  DFFSRHQX4TS addWeight_7__add_S_reg_0_ ( .D(addWeight_7__add_s[0]), .CK(clk), 
        .SN(n79), .RN(n80), .Q(n2430) );
  DFFSRHQX4TS addWeight_13__add_S_reg_0_ ( .D(addWeight_13__add_s[0]), .CK(clk), .SN(n139), .RN(n140), .Q(n2413) );
  DFFSRHQX4TS addWeight_14__add_S_reg_0_ ( .D(addWeight_14__add_s[0]), .CK(clk), .SN(n149), .RN(n150), .Q(n2410) );
  DFFSRHQX4TS addWeight_18__add_S_reg_0_ ( .D(addWeight_18__add_s[0]), .CK(clk), .SN(n189), .RN(n190), .Q(n2399) );
  DFFSRHQX4TS addWeight_4__add_S_reg_0_ ( .D(addWeight_4__add_s[0]), .CK(clk), 
        .SN(n49), .RN(n50), .Q(n2439) );
  DFFSRHQX4TS addWeight_5__add_S_reg_0_ ( .D(addWeight_5__add_s[0]), .CK(clk), 
        .SN(n59), .RN(n60), .Q(n2436) );
  DFFSRHQX4TS addWeight_3__add_S_reg_0_ ( .D(addWeight_3__add_s[0]), .CK(clk), 
        .SN(n39), .RN(n40), .Q(n2442) );
  DFFSRHQX4TS addWeight_16__add_S_reg_0_ ( .D(addWeight_16__add_s[0]), .CK(clk), .SN(n169), .RN(n170), .Q(sumOut[128]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_1_ ( .D(addWeight_2__add_s[1]), .CK(clk), 
        .SN(n21), .RN(n22), .Q(sumOut[17]) );
  DFFSRHQX4TS addWeight_12__add_S_reg_0_ ( .D(addWeight_12__add_s[0]), .CK(clk), .SN(n129), .RN(n130), .Q(n2416) );
  DFFSRHQX4TS addWeight_28__add_S_reg_0_ ( .D(addWeight_28__add_s[0]), .CK(clk), .SN(n289), .RN(n290), .Q(sumOut[224]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_0_ ( .D(addWeight_11__add_s[0]), .CK(clk), .SN(n119), .RN(n120), .Q(n2419) );
  DFFSRHQX4TS addWeight_1__add_S_reg_0_ ( .D(addWeight_1__add_s[0]), .CK(clk), 
        .SN(n19), .RN(n20), .Q(n2446) );
  DFFSRHQX4TS addWeight_6__add_S_reg_4_ ( .D(addWeight_6__add_s[4]), .CK(clk), 
        .SN(n67), .RN(n68), .Q(sumOut[52]) );
  DFFSRHQX4TS addWeight_19__add_S_reg_4_ ( .D(addWeight_19__add_s[4]), .CK(clk), .SN(n197), .RN(n198), .Q(sumOut[156]) );
  DFFSRHQX4TS addWeight_20__add_S_reg_4_ ( .D(addWeight_20__add_s[4]), .CK(clk), .SN(n207), .RN(n208), .Q(sumOut[164]) );
  DFFSRHQX4TS addWeight_30__add_S_reg_4_ ( .D(addWeight_30__add_s[4]), .CK(clk), .SN(n307), .RN(n308), .Q(sumOut[244]) );
  DFFSRHQX4TS addWeight_23__add_S_reg_4_ ( .D(addWeight_23__add_s[4]), .CK(clk), .SN(n237), .RN(n238), .Q(sumOut[188]) );
  DFFSRHQX4TS addWeight_24__add_S_reg_4_ ( .D(addWeight_24__add_s[4]), .CK(clk), .SN(n247), .RN(n248), .Q(sumOut[196]) );
  DFFSRHQX4TS addWeight_22__add_S_reg_4_ ( .D(addWeight_22__add_s[4]), .CK(clk), .SN(n227), .RN(n228), .Q(sumOut[180]) );
  DFFSRHQX4TS addWeight_4__add_S_reg_4_ ( .D(addWeight_4__add_s[4]), .CK(clk), 
        .SN(n47), .RN(n48), .Q(sumOut[36]) );
  DFFSRHQX4TS addWeight_5__add_S_reg_4_ ( .D(addWeight_5__add_s[4]), .CK(clk), 
        .SN(n57), .RN(n58), .Q(sumOut[44]) );
  DFFSRHQX4TS addWeight_3__add_S_reg_4_ ( .D(addWeight_3__add_s[4]), .CK(clk), 
        .SN(n37), .RN(n38), .Q(sumOut[28]) );
  DFFSRHQX4TS addWeight_26__add_S_reg_4_ ( .D(addWeight_26__add_s[4]), .CK(clk), .SN(n267), .RN(n268), .Q(sumOut[212]) );
  DFFSRHQX4TS addWeight_21__add_S_reg_4_ ( .D(addWeight_21__add_s[4]), .CK(clk), .SN(n217), .RN(n218), .Q(sumOut[172]) );
  DFFSRHQX4TS addWeight_12__add_S_reg_4_ ( .D(addWeight_12__add_s[4]), .CK(clk), .SN(n127), .RN(n128), .Q(sumOut[100]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_4_ ( .D(addWeight_29__add_s[4]), .CK(clk), .SN(n297), .RN(n298), .Q(sumOut[236]) );
  DFFSRHQX4TS addWeight_31__add_S_reg_4_ ( .D(addWeight_31__add_s[4]), .CK(clk), .SN(n317), .RN(n318), .Q(sumOut[252]) );
  DFFSRHQX4TS addWeight_10__add_S_reg_4_ ( .D(addWeight_10__add_s[4]), .CK(clk), .SN(n107), .RN(n108), .Q(sumOut[84]) );
  DFFSRHQX4TS addWeight_0__add_S_reg_4_ ( .D(addWeight_0__add_s[4]), .CK(clk), 
        .SN(n7), .RN(n8), .Q(sumOut[4]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_4_ ( .D(addWeight_11__add_s[4]), .CK(clk), .SN(n117), .RN(n118), .Q(sumOut[92]) );
  DFFSRHQX4TS addWeight_1__add_S_reg_4_ ( .D(addWeight_1__add_s[4]), .CK(clk), 
        .SN(n17), .RN(n18), .Q(sumOut[12]) );
  DFFSRHQX4TS addWeight_28__add_S_reg_4_ ( .D(addWeight_28__add_s[4]), .CK(clk), .SN(n287), .RN(n288), .Q(sumOut[228]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_0_ ( .D(addWeight_2__add_s[0]), .CK(clk), 
        .SN(n29), .RN(n30), .Q(sumOut[16]) );
  DFFSRHQX4TS addWeight_26__add_S_reg_2_ ( .D(addWeight_26__add_s[2]), .CK(clk), .SN(n263), .RN(n264), .Q(sumOut[210]) );
  DFFSRHQX4TS addWeight_12__add_S_reg_5_ ( .D(addWeight_12__add_s[5]), .CK(clk), .SN(n127), .RN(n128), .Q(sumOut[101]) );
  DFFSRHQX4TS addWeight_27__add_S_reg_6_ ( .D(addWeight_27__add_s[6]), .CK(clk), .SN(n277), .RN(n278), .Q(sumOut[222]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_6_ ( .D(addWeight_2__add_s[6]), .CK(clk), 
        .SN(n27), .RN(n28), .Q(sumOut[22]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_7_ ( .D(addWeight_2__add_s[7]), .CK(clk), 
        .SN(n27), .RN(n28), .Q(sumOut[23]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_4_ ( .D(addWeight_2__add_s[4]), .CK(clk), 
        .SN(n27), .RN(n28), .Q(sumOut[20]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_5_ ( .D(addWeight_29__add_s[5]), .CK(clk), .SN(n297), .RN(n298), .Q(sumOut[237]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_5_ ( .D(addWeight_11__add_s[5]), .CK(clk), .SN(n117), .RN(n118), .Q(sumOut[93]) );
  DFFSRHQX4TS addWeight_1__add_S_reg_5_ ( .D(addWeight_1__add_s[5]), .CK(clk), 
        .SN(n17), .RN(n18), .Q(sumOut[13]) );
  DFFSRHQX4TS addWeight_27__add_S_reg_7_ ( .D(addWeight_27__add_s[7]), .CK(clk), .SN(n277), .RN(n278), .Q(sumOut[223]) );
  DFFSRHQX4TS addWeight_10__add_S_reg_5_ ( .D(addWeight_10__add_s[5]), .CK(clk), .SN(n107), .RN(n108), .Q(sumOut[85]) );
  DFFSRHQX4TS addWeight_12__add_S_reg_6_ ( .D(addWeight_12__add_s[6]), .CK(clk), .SN(n127), .RN(n128), .Q(sumOut[102]) );
  DFFSRHQX4TS addWeight_0__add_S_reg_5_ ( .D(addWeight_0__add_s[5]), .CK(clk), 
        .SN(n7), .RN(n8), .Q(sumOut[5]) );
  DFFSRHQX4TS addWeight_31__add_S_reg_5_ ( .D(addWeight_31__add_s[5]), .CK(clk), .SN(n317), .RN(n318), .Q(sumOut[253]) );
  DFFSRHQX4TS addWeight_12__add_S_reg_7_ ( .D(addWeight_12__add_s[7]), .CK(clk), .SN(n127), .RN(n128), .Q(sumOut[103]) );
  DFFSRHQX4TS addWeight_26__add_S_reg_5_ ( .D(addWeight_26__add_s[5]), .CK(clk), .SN(n267), .RN(n268), .Q(sumOut[213]) );
  DFFSRHQX4TS addWeight_2__add_S_reg_3_ ( .D(addWeight_2__add_s[3]), .CK(clk), 
        .SN(n25), .RN(n26), .Q(n2443) );
  DFFSRHQX4TS addWeight_25__add_S_reg_7_ ( .D(addWeight_25__add_s[7]), .CK(clk), .SN(n257), .RN(n258), .Q(sumOut[207]) );
  DFFSRHQX4TS addWeight_16__add_S_reg_5_ ( .D(addWeight_16__add_s[5]), .CK(clk), .SN(n167), .RN(n168), .Q(sumOut[133]) );
  DFFSRHQX4TS addWeight_15__add_S_reg_5_ ( .D(addWeight_15__add_s[5]), .CK(clk), .SN(n157), .RN(n158), .Q(sumOut[125]) );
  DFFSRHQX4TS addWeight_7__add_S_reg_5_ ( .D(addWeight_7__add_s[5]), .CK(clk), 
        .SN(n77), .RN(n78), .Q(sumOut[61]) );
  DFFSRHQX4TS addWeight_6__add_S_reg_5_ ( .D(addWeight_6__add_s[5]), .CK(clk), 
        .SN(n67), .RN(n68), .Q(sumOut[53]) );
  DFFSRHQX4TS addWeight_5__add_S_reg_5_ ( .D(addWeight_5__add_s[5]), .CK(clk), 
        .SN(n57), .RN(n58), .Q(sumOut[45]) );
  DFFSRHQX4TS addWeight_4__add_S_reg_5_ ( .D(addWeight_4__add_s[5]), .CK(clk), 
        .SN(n47), .RN(n48), .Q(sumOut[37]) );
  DFFSRHQX4TS addWeight_3__add_S_reg_5_ ( .D(addWeight_3__add_s[5]), .CK(clk), 
        .SN(n37), .RN(n38), .Q(sumOut[29]) );
  DFFSRHQX4TS addWeight_18__add_S_reg_5_ ( .D(addWeight_18__add_s[5]), .CK(clk), .SN(n187), .RN(n188), .Q(sumOut[149]) );
  DFFSRHQX4TS addWeight_17__add_S_reg_5_ ( .D(addWeight_17__add_s[5]), .CK(clk), .SN(n177), .RN(n178), .Q(sumOut[141]) );
  DFFSRHQX4TS addWeight_14__add_S_reg_5_ ( .D(addWeight_14__add_s[5]), .CK(clk), .SN(n147), .RN(n148), .Q(sumOut[117]) );
  DFFSRHQX4TS addWeight_13__add_S_reg_5_ ( .D(addWeight_13__add_s[5]), .CK(clk), .SN(n137), .RN(n138), .Q(sumOut[109]) );
  DFFSRHQX4TS addWeight_9__add_S_reg_5_ ( .D(addWeight_9__add_s[5]), .CK(clk), 
        .SN(n97), .RN(n98), .Q(sumOut[77]) );
  DFFSRHQX4TS addWeight_8__add_S_reg_5_ ( .D(addWeight_8__add_s[5]), .CK(clk), 
        .SN(n87), .RN(n88), .Q(sumOut[69]) );
  DFFSRHQX4TS addWeight_28__add_S_reg_5_ ( .D(addWeight_28__add_s[5]), .CK(clk), .SN(n287), .RN(n288), .Q(sumOut[229]) );
  DFFSRHQX4TS addWeight_26__add_S_reg_6_ ( .D(addWeight_26__add_s[6]), .CK(clk), .SN(n267), .RN(n268), .Q(sumOut[214]) );
  DFFSRHQX4TS addWeight_10__add_S_reg_7_ ( .D(addWeight_10__add_s[7]), .CK(clk), .SN(n107), .RN(n108), .Q(sumOut[87]) );
  DFFSRHQX4TS addWeight_28__add_S_reg_7_ ( .D(addWeight_28__add_s[7]), .CK(clk), .SN(n287), .RN(n288), .Q(sumOut[231]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_6_ ( .D(addWeight_29__add_s[6]), .CK(clk), .SN(n297), .RN(n298), .Q(sumOut[238]) );
  DFFSRHQX4TS addWeight_29__add_S_reg_7_ ( .D(addWeight_29__add_s[7]), .CK(clk), .SN(n297), .RN(n298), .Q(sumOut[239]) );
  DFFSRHQX4TS addWeight_27__add_S_reg_4_ ( .D(addWeight_27__add_s[4]), .CK(clk), .SN(n277), .RN(n278), .Q(sumOut[220]) );
  DFFSRHQX4TS addWeight_27__add_S_reg_3_ ( .D(addWeight_27__add_s[3]), .CK(clk), .SN(n275), .RN(n276), .Q(n2378) );
  DFFSRHQX4TS addWeight_18__add_S_reg_6_ ( .D(addWeight_18__add_s[6]), .CK(clk), .SN(n187), .RN(n188), .Q(sumOut[150]) );
  DFFSRHQX4TS addWeight_17__add_S_reg_6_ ( .D(addWeight_17__add_s[6]), .CK(clk), .SN(n177), .RN(n178), .Q(sumOut[142]) );
  DFFSRHQX4TS addWeight_16__add_S_reg_6_ ( .D(addWeight_16__add_s[6]), .CK(clk), .SN(n167), .RN(n168), .Q(sumOut[134]) );
  DFFSRHQX4TS addWeight_15__add_S_reg_6_ ( .D(addWeight_15__add_s[6]), .CK(clk), .SN(n157), .RN(n158), .Q(sumOut[126]) );
  DFFSRHQX4TS addWeight_14__add_S_reg_6_ ( .D(addWeight_14__add_s[6]), .CK(clk), .SN(n147), .RN(n148), .Q(sumOut[118]) );
  DFFSRHQX4TS addWeight_13__add_S_reg_6_ ( .D(addWeight_13__add_s[6]), .CK(clk), .SN(n137), .RN(n138), .Q(sumOut[110]) );
  DFFSRHQX4TS addWeight_9__add_S_reg_6_ ( .D(addWeight_9__add_s[6]), .CK(clk), 
        .SN(n97), .RN(n98), .Q(sumOut[78]) );
  DFFSRHQX4TS addWeight_8__add_S_reg_6_ ( .D(addWeight_8__add_s[6]), .CK(clk), 
        .SN(n87), .RN(n88), .Q(sumOut[70]) );
  DFFSRHQX4TS addWeight_7__add_S_reg_6_ ( .D(addWeight_7__add_s[6]), .CK(clk), 
        .SN(n77), .RN(n78), .Q(sumOut[62]) );
  DFFSRHQX4TS addWeight_6__add_S_reg_6_ ( .D(addWeight_6__add_s[6]), .CK(clk), 
        .SN(n67), .RN(n68), .Q(sumOut[54]) );
  DFFSRHQX4TS addWeight_5__add_S_reg_6_ ( .D(addWeight_5__add_s[6]), .CK(clk), 
        .SN(n57), .RN(n58), .Q(sumOut[46]) );
  DFFSRHQX4TS addWeight_4__add_S_reg_6_ ( .D(addWeight_4__add_s[6]), .CK(clk), 
        .SN(n47), .RN(n48), .Q(sumOut[38]) );
  DFFSRHQX4TS addWeight_3__add_S_reg_6_ ( .D(addWeight_3__add_s[6]), .CK(clk), 
        .SN(n37), .RN(n38), .Q(sumOut[30]) );
  DFFSRHQX4TS addWeight_26__add_S_reg_7_ ( .D(addWeight_26__add_s[7]), .CK(clk), .SN(n267), .RN(n268), .Q(sumOut[215]) );
  DFFSRHQX4TS addWeight_26__add_S_reg_3_ ( .D(addWeight_26__add_s[3]), .CK(clk), .SN(n265), .RN(n266), .Q(n2379) );
  DFFSRHQX4TS addWeight_18__add_S_reg_4_ ( .D(addWeight_18__add_s[4]), .CK(clk), .SN(n187), .RN(n188), .Q(sumOut[148]) );
  DFFSRHQX4TS addWeight_17__add_S_reg_4_ ( .D(addWeight_17__add_s[4]), .CK(clk), .SN(n177), .RN(n178), .Q(sumOut[140]) );
  DFFSRHQX4TS addWeight_16__add_S_reg_4_ ( .D(addWeight_16__add_s[4]), .CK(clk), .SN(n167), .RN(n168), .Q(sumOut[132]) );
  DFFSRHQX4TS addWeight_15__add_S_reg_4_ ( .D(addWeight_15__add_s[4]), .CK(clk), .SN(n157), .RN(n158), .Q(sumOut[124]) );
  DFFSRHQX4TS addWeight_14__add_S_reg_4_ ( .D(addWeight_14__add_s[4]), .CK(clk), .SN(n147), .RN(n148), .Q(sumOut[116]) );
  DFFSRHQX4TS addWeight_13__add_S_reg_4_ ( .D(addWeight_13__add_s[4]), .CK(clk), .SN(n137), .RN(n138), .Q(sumOut[108]) );
  DFFSRHQX4TS addWeight_9__add_S_reg_4_ ( .D(addWeight_9__add_s[4]), .CK(clk), 
        .SN(n97), .RN(n98), .Q(sumOut[76]) );
  DFFSRHQX4TS addWeight_8__add_S_reg_4_ ( .D(addWeight_8__add_s[4]), .CK(clk), 
        .SN(n87), .RN(n88), .Q(sumOut[68]) );
  DFFSRHQX4TS addWeight_7__add_S_reg_4_ ( .D(addWeight_7__add_s[4]), .CK(clk), 
        .SN(n77), .RN(n78), .Q(sumOut[60]) );
  DFFSRHQX4TS addWeight_19__add_S_reg_0_ ( .D(addWeight_19__add_s[0]), .CK(clk), .SN(n199), .RN(n200), .Q(sumOut[152]) );
  DFFSRHQX4TS addWeight_20__add_S_reg_0_ ( .D(addWeight_20__add_s[0]), .CK(clk), .SN(n209), .RN(n210), .Q(n2394) );
  DFFSRHQX4TS addWeight_23__add_S_reg_0_ ( .D(addWeight_23__add_s[0]), .CK(clk), .SN(n239), .RN(n240), .Q(sumOut[184]) );
  DFFSRHQX4TS addWeight_24__add_S_reg_0_ ( .D(addWeight_24__add_s[0]), .CK(clk), .SN(n249), .RN(n250), .Q(n2385) );
  DFFSRHQX4TS addWeight_21__add_S_reg_0_ ( .D(addWeight_21__add_s[0]), .CK(clk), .SN(n219), .RN(n220), .Q(sumOut[168]) );
  DFFSRHQX4TS addWeight_22__add_S_reg_0_ ( .D(addWeight_22__add_s[0]), .CK(clk), .SN(n229), .RN(n230), .Q(sumOut[176]) );
  DFFSRHQX4TS addWeight_30__add_S_reg_0_ ( .D(addWeight_30__add_s[0]), .CK(clk), .SN(n309), .RN(n310), .Q(sumOut[240]) );
  DFFSRHQX4TS addWeight_31__add_S_reg_6_ ( .D(addWeight_31__add_s[6]), .CK(clk), .SN(n317), .RN(n318), .Q(sumOut[254]) );
  DFFSRHQX4TS addWeight_0__add_S_reg_6_ ( .D(addWeight_0__add_s[6]), .CK(clk), 
        .SN(n7), .RN(n8), .Q(sumOut[6]) );
  DFFSRHQX4TS addWeight_11__add_S_reg_6_ ( .D(addWeight_11__add_s[6]), .CK(clk), .SN(n117), .RN(n118), .Q(sumOut[94]) );
  DFFSRHQX4TS addWeight_10__add_S_reg_6_ ( .D(addWeight_10__add_s[6]), .CK(clk), .SN(n107), .RN(n108), .Q(sumOut[86]) );
  DFFSRHQX4TS addWeight_19__add_S_reg_6_ ( .D(addWeight_19__add_s[6]), .CK(clk), .SN(n197), .RN(n198), .Q(sumOut[158]) );
  DFFSRHQX4TS addWeight_28__add_S_reg_6_ ( .D(addWeight_28__add_s[6]), .CK(clk), .SN(n287), .RN(n288), .Q(sumOut[230]) );
  AOI2BB1X1TS U322 ( .A0N(sumOut[248]), .A1N(n556), .B0(n715), .Y(
        addWeight_31__add_s[0]) );
  XOR2X1TS U323 ( .A(n542), .B(n762), .Y(addWeight_28__add_s[3]) );
  CLKBUFX2TS U324 ( .A(n2374), .Y(sumOut[234]) );
  CLKBUFX2TS U325 ( .A(n2443), .Y(sumOut[19]) );
  CLKBUFX2TS U326 ( .A(n2396), .Y(sumOut[154]) );
  CLKBUFX2TS U327 ( .A(n2421), .Y(sumOut[82]) );
  OAI2BB1X2TS U328 ( .A0N(n1411), .A1N(n1790), .B0(n1410), .Y(n1415) );
  NAND2X1TS U329 ( .A(n2235), .B(n2234), .Y(n2236) );
  NAND2X1TS U330 ( .A(n727), .B(n728), .Y(n729) );
  NAND2X1TS U331 ( .A(n712), .B(n1524), .Y(n713) );
  NAND2X1TS U332 ( .A(n625), .B(n624), .Y(n626) );
  NAND2XLTS U333 ( .A(n769), .B(n768), .Y(n770) );
  NAND2XLTS U334 ( .A(n744), .B(n1447), .Y(n745) );
  NAND2XLTS U335 ( .A(n778), .B(n777), .Y(n779) );
  NOR2X1TS U336 ( .A(n1557), .B(n1556), .Y(n616) );
  NAND2BX2TS U337 ( .AN(n466), .B(n1426), .Y(n1431) );
  INVX4TS U338 ( .A(n1537), .Y(n322) );
  CLKAND2X2TS U339 ( .A(n1105), .B(n1103), .Y(n866) );
  NOR2XLTS U340 ( .A(n1548), .B(n1547), .Y(n655) );
  NOR2XLTS U341 ( .A(n1539), .B(n1538), .Y(n663) );
  NAND2X1TS U342 ( .A(n1499), .B(n1498), .Y(n357) );
  AND2X2TS U343 ( .A(n1175), .B(n1173), .Y(n951) );
  NAND2X1TS U344 ( .A(n749), .B(n1459), .Y(n1639) );
  NAND2X1TS U345 ( .A(n1856), .B(n1855), .Y(n2249) );
  NAND2X1TS U346 ( .A(n1997), .B(n1996), .Y(n2224) );
  NAND2X1TS U347 ( .A(n1893), .B(n1892), .Y(n2219) );
  NAND2X1TS U348 ( .A(n1838), .B(n1837), .Y(n2184) );
  NAND2X1TS U349 ( .A(n1978), .B(n1977), .Y(n2174) );
  NAND2XLTS U350 ( .A(n1496), .B(n1499), .Y(n464) );
  NOR2X1TS U351 ( .A(n1249), .B(n1813), .Y(n1256) );
  NOR2X1TS U352 ( .A(n1388), .B(n1744), .Y(n1086) );
  NOR2X1TS U353 ( .A(n1370), .B(n1764), .Y(n1116) );
  NOR2X1TS U354 ( .A(n1376), .B(n1726), .Y(n1106) );
  NOR2X1TS U355 ( .A(n1340), .B(n1773), .Y(n1166) );
  NOR2X1TS U356 ( .A(n1364), .B(n1778), .Y(n1126) );
  NOR2X1TS U357 ( .A(n1358), .B(n1759), .Y(n1136) );
  NOR2X1TS U358 ( .A(n1328), .B(n1783), .Y(n1186) );
  NOR2X1TS U359 ( .A(n1412), .B(n1787), .Y(n1046) );
  NOR2X1TS U360 ( .A(n1400), .B(n1800), .Y(n1066) );
  NOR2X1TS U361 ( .A(n1394), .B(n1804), .Y(n1076) );
  NOR2X1TS U362 ( .A(n1316), .B(n1749), .Y(n1206) );
  NOR2X1TS U363 ( .A(n1322), .B(n1731), .Y(n1196) );
  NOR2BX2TS U364 ( .AN(n1281), .B(n578), .Y(n581) );
  NOR2X1TS U365 ( .A(n1561), .B(n1557), .Y(n1478) );
  OR2X2TS U366 ( .A(sumOut[202]), .B(n725), .Y(n2234) );
  NAND2BX1TS U367 ( .AN(n1473), .B(sumOut[102]), .Y(n1504) );
  NOR2BX2TS U368 ( .AN(n601), .B(n618), .Y(n642) );
  AOI21X2TS U369 ( .A0(sumOut[207]), .A1(n1536), .B0(n1535), .Y(n1537) );
  NAND2X2TS U370 ( .A(n1565), .B(n1568), .Y(n548) );
  NOR2X2TS U371 ( .A(n1286), .B(n2012), .Y(n1273) );
  NAND2BX1TS U372 ( .AN(n1527), .B(sumOut[6]), .Y(n1574) );
  NAND2BXLTS U373 ( .AN(n582), .B(sumOut[86]), .Y(n1282) );
  INVX2TS U374 ( .A(n1280), .Y(n578) );
  CLKAND2X2TS U375 ( .A(sumOut[236]), .B(n1270), .Y(n1808) );
  NAND2BX1TS U376 ( .AN(sumOut[102]), .B(n1473), .Y(n1503) );
  NOR2X1TS U377 ( .A(n2011), .B(n1287), .Y(n1274) );
  NOR2X2TS U378 ( .A(n1579), .B(n2024), .Y(n1571) );
  INVX4TS U379 ( .A(n532), .Y(n531) );
  INVX4TS U380 ( .A(n520), .Y(n519) );
  NAND2BX2TS U381 ( .AN(n480), .B(n1572), .Y(n479) );
  NAND2BX2TS U382 ( .AN(sumOut[230]), .B(n1435), .Y(n1480) );
  NAND2X2TS U383 ( .A(n2141), .B(n1649), .Y(n701) );
  CLKINVX3TS U384 ( .A(n1603), .Y(n764) );
  NOR2X1TS U385 ( .A(n1547), .B(n1553), .Y(n1485) );
  NAND2X1TS U386 ( .A(n595), .B(n594), .Y(n644) );
  NOR2X1TS U387 ( .A(sumOut[21]), .B(n1260), .Y(n1248) );
  NOR2X1TS U388 ( .A(sumOut[245]), .B(n1050), .Y(n1413) );
  NOR2X1TS U389 ( .A(sumOut[197]), .B(n1060), .Y(n1407) );
  NOR2X1TS U390 ( .A(sumOut[189]), .B(n1070), .Y(n1401) );
  NOR2X1TS U391 ( .A(sumOut[181]), .B(n1080), .Y(n1395) );
  NOR2X1TS U392 ( .A(sumOut[173]), .B(n1090), .Y(n1389) );
  NOR2X1TS U393 ( .A(sumOut[165]), .B(n1100), .Y(n1383) );
  NOR2X1TS U394 ( .A(sumOut[157]), .B(n1110), .Y(n1377) );
  NOR2X1TS U395 ( .A(sumOut[149]), .B(n1120), .Y(n1371) );
  NOR2X1TS U396 ( .A(sumOut[133]), .B(n1140), .Y(n1359) );
  NOR2X1TS U397 ( .A(sumOut[125]), .B(n1150), .Y(n1353) );
  NOR2X1TS U398 ( .A(sumOut[117]), .B(n1160), .Y(n1347) );
  NOR2X1TS U399 ( .A(sumOut[109]), .B(n1170), .Y(n1341) );
  NOR2X1TS U400 ( .A(sumOut[77]), .B(n1180), .Y(n1335) );
  NOR2X1TS U401 ( .A(sumOut[69]), .B(n1190), .Y(n1329) );
  NOR2X1TS U402 ( .A(sumOut[61]), .B(n1200), .Y(n1323) );
  NOR2X1TS U403 ( .A(sumOut[53]), .B(n1210), .Y(n1317) );
  NOR2X1TS U404 ( .A(sumOut[45]), .B(n1220), .Y(n1311) );
  NOR2X1TS U405 ( .A(sumOut[37]), .B(n1230), .Y(n1305) );
  NOR2X1TS U406 ( .A(sumOut[29]), .B(n1240), .Y(n1299) );
  NOR2X1TS U407 ( .A(sumOut[237]), .B(n1270), .Y(n1243) );
  NOR2X1TS U408 ( .A(sumOut[213]), .B(n1456), .Y(n1515) );
  NOR2X2TS U409 ( .A(n700), .B(n568), .Y(n2141) );
  NOR2X2TS U410 ( .A(sumOut[228]), .B(n1437), .Y(n1556) );
  NOR2X2TS U411 ( .A(sumOut[252]), .B(n1040), .Y(n2011) );
  NOR2X2TS U412 ( .A(sumOut[12]), .B(n1421), .Y(n1538) );
  NAND2X2TS U413 ( .A(n1029), .B(n1667), .Y(n1033) );
  NAND2X2TS U414 ( .A(n1518), .B(n1521), .Y(n475) );
  NOR2X2TS U415 ( .A(n617), .B(n593), .Y(n643) );
  NOR2X2TS U416 ( .A(n2019), .B(n1293), .Y(n1280) );
  AND2X6TS U417 ( .A(sumOut[203]), .B(n664), .Y(n726) );
  AND2X6TS U418 ( .A(sumOut[218]), .B(n559), .Y(n2263) );
  OR2X6TS U419 ( .A(n2435), .B(n401), .Y(n532) );
  OR2X6TS U420 ( .A(n2409), .B(n414), .Y(n520) );
  BUFX3TS U421 ( .A(n2414), .Y(sumOut[99]) );
  INVX2TS U422 ( .A(n1416), .Y(n1421) );
  INVX6TS U423 ( .A(n332), .Y(n1614) );
  INVX2TS U424 ( .A(n1035), .Y(n1040) );
  OR2X4TS U425 ( .A(n2415), .B(n1463), .Y(n1599) );
  NOR2X2TS U426 ( .A(sumOut[4]), .B(n1529), .Y(n2023) );
  AND2X4TS U427 ( .A(sumOut[2]), .B(n710), .Y(n1618) );
  AND2X4TS U428 ( .A(sumOut[210]), .B(n1440), .Y(n1628) );
  OR2X4TS U429 ( .A(n2372), .B(n1709), .Y(n1936) );
  OR2X4TS U430 ( .A(n2384), .B(n1654), .Y(n1946) );
  OR2X4TS U431 ( .A(n2387), .B(n1704), .Y(n1956) );
  OR2X4TS U432 ( .A(n2389), .B(n1691), .Y(n1966) );
  OR2X4TS U433 ( .A(n2391), .B(n1663), .Y(n1985) );
  OR2X4TS U434 ( .A(n2393), .B(n1673), .Y(n1881) );
  INVX2TS U435 ( .A(n1432), .Y(n1437) );
  AND2X4TS U436 ( .A(n2380), .B(n725), .Y(n2233) );
  INVX2TS U437 ( .A(n932), .Y(n933) );
  INVX2TS U438 ( .A(n897), .Y(n898) );
  INVX2TS U439 ( .A(n969), .Y(n970) );
  INVX2TS U440 ( .A(n799), .Y(n800) );
  INVX2TS U441 ( .A(n849), .Y(n850) );
  INVX2TS U442 ( .A(n1006), .Y(n1007) );
  INVX2TS U443 ( .A(n945), .Y(n946) );
  INVX2TS U444 ( .A(n711), .Y(n1519) );
  CLKBUFX2TS U445 ( .A(weightsIn[96]), .Y(n1682) );
  INVX2TS U446 ( .A(n363), .Y(n364) );
  INVX2TS U447 ( .A(n664), .Y(n323) );
  CLKBUFX2TS U448 ( .A(weightsIn[145]), .Y(n2172) );
  CLKBUFX2TS U449 ( .A(weightsIn[50]), .Y(n2142) );
  CLKBUFX2TS U450 ( .A(weightsIn[2]), .Y(n710) );
  CLKBUFX2TS U451 ( .A(weightsIn[137]), .Y(n559) );
  INVX2TS U452 ( .A(n1424), .Y(n1429) );
  CLKBUFX2TS U453 ( .A(weightsIn[77]), .Y(n905) );
  CLKBUFX2TS U454 ( .A(weightsIn[72]), .Y(n917) );
  CLKBUFX2TS U455 ( .A(weightsIn[92]), .Y(n869) );
  CLKBUFX2TS U456 ( .A(weightsIn[17]), .Y(n1015) );
  CLKBUFX2TS U457 ( .A(weightsIn[27]), .Y(n990) );
  CLKBUFX2TS U458 ( .A(weightsIn[62]), .Y(n750) );
  CLKBUFX2TS U459 ( .A(weightsIn[142]), .Y(n612) );
  CLKBUFX2TS U460 ( .A(weightsIn[57]), .Y(n651) );
  CLKBUFX2TS U461 ( .A(weightsIn[7]), .Y(n659) );
  INVX2TS U462 ( .A(n564), .Y(n605) );
  INVX1TS U463 ( .A(n1019), .Y(n337) );
  INVX1TS U464 ( .A(n873), .Y(n338) );
  INVX1TS U465 ( .A(n994), .Y(n339) );
  INVX1TS U466 ( .A(n921), .Y(n340) );
  INVX1TS U467 ( .A(n826), .Y(n341) );
  INVX1TS U468 ( .A(n813), .Y(n342) );
  INVX1TS U469 ( .A(n787), .Y(n343) );
  INVX1TS U470 ( .A(n982), .Y(n344) );
  INVX1TS U471 ( .A(n909), .Y(n345) );
  INVX1TS U472 ( .A(n886), .Y(n346) );
  INVX1TS U473 ( .A(n958), .Y(n347) );
  BUFX3TS U474 ( .A(weightsIn[128]), .Y(n664) );
  BUFX2TS U475 ( .A(weightsIn[158]), .Y(n1026) );
  BUFX2TS U476 ( .A(weightsIn[63]), .Y(n751) );
  BUFX2TS U477 ( .A(weightsIn[148]), .Y(n678) );
  INVX2TS U478 ( .A(n361), .Y(n362) );
  CLKINVX2TS U479 ( .A(n884), .Y(n485) );
  CLKINVX2TS U480 ( .A(n944), .Y(n500) );
  CLKINVX2TS U481 ( .A(n1005), .Y(n511) );
  INVX2TS U482 ( .A(n371), .Y(n372) );
  INVX2TS U483 ( .A(n373), .Y(n374) );
  CLKBUFX2TS U484 ( .A(weightsIn[140]), .Y(n2164) );
  INVX2TS U485 ( .A(weightsIn[23]), .Y(n1006) );
  INVX2TS U486 ( .A(weightsIn[48]), .Y(n945) );
  INVX2TS U487 ( .A(weightsIn[68]), .Y(n932) );
  INVX2TS U488 ( .A(weightsIn[83]), .Y(n897) );
  INVX2TS U489 ( .A(weightsIn[103]), .Y(n849) );
  INVX2TS U490 ( .A(weightsIn[123]), .Y(n799) );
  INVX2TS U491 ( .A(weightsIn[38]), .Y(n969) );
  CLKBUFX2TS U492 ( .A(weightsIn[125]), .Y(n2146) );
  INVX2TS U493 ( .A(weightsIn[13]), .Y(n686) );
  INVX2TS U494 ( .A(n1525), .Y(n1526) );
  BUFX3TS U495 ( .A(weightsIn[15]), .Y(n1017) );
  BUFX3TS U496 ( .A(weightsIn[25]), .Y(n992) );
  BUFX3TS U497 ( .A(weightsIn[90]), .Y(n871) );
  BUFX3TS U498 ( .A(weightsIn[70]), .Y(n919) );
  BUFX3TS U499 ( .A(weightsIn[65]), .Y(n931) );
  BUFX3TS U500 ( .A(weightsIn[35]), .Y(n968) );
  BUFX3TS U501 ( .A(weightsIn[75]), .Y(n907) );
  BUFX3TS U502 ( .A(weightsIn[30]), .Y(n980) );
  BUFX3TS U503 ( .A(weightsIn[40]), .Y(n956) );
  CLKBUFX2TS U504 ( .A(weightsIn[0]), .Y(n2153) );
  CLKBUFX2TS U505 ( .A(weightsIn[133]), .Y(n743) );
  CLKINVX2TS U506 ( .A(n400), .Y(n402) );
  CLKINVX2TS U507 ( .A(n417), .Y(n419) );
  CLKBUFX2TS U508 ( .A(weightsIn[55]), .Y(n2167) );
  CLKBUFX2TS U509 ( .A(weightsIn[5]), .Y(n2170) );
  CLKBUFX2TS U510 ( .A(weightsIn[155]), .Y(n556) );
  CLKBUFX2TS U511 ( .A(weightsIn[80]), .Y(n896) );
  INVX2TS U512 ( .A(n413), .Y(n414) );
  CLKINVX2TS U513 ( .A(weightsIn[8]), .Y(n375) );
  CLKINVX2TS U514 ( .A(weightsIn[58]), .Y(n379) );
  CLKINVX2TS U515 ( .A(weightsIn[108]), .Y(n387) );
  CLKINVX2TS U516 ( .A(weightsIn[143]), .Y(n391) );
  AOI21X1TS U517 ( .A0(n2177), .A1(n2174), .B0(n2173), .Y(n1983) );
  AOI21X1TS U518 ( .A0(n2227), .A1(n2224), .B0(n2223), .Y(n2002) );
  BUFX4TS U519 ( .A(n2373), .Y(sumOut[235]) );
  BUFX4TS U520 ( .A(n2404), .Y(sumOut[129]) );
  OAI21X2TS U521 ( .A0(n1976), .A1(n535), .B0(n1975), .Y(n2177) );
  CLKINVX3TS U522 ( .A(n536), .Y(n535) );
  OAI21X2TS U523 ( .A0(n1995), .A1(n517), .B0(n1994), .Y(n2227) );
  CLKINVX3TS U524 ( .A(n518), .Y(n517) );
  NAND2X2TS U525 ( .A(n2441), .B(n372), .Y(n513) );
  BUFX4TS U526 ( .A(n2441), .Y(sumOut[25]) );
  NAND2X2TS U527 ( .A(n2406), .B(n374), .Y(n493) );
  BUFX4TS U528 ( .A(n2406), .Y(sumOut[121]) );
  AND2X4TS U529 ( .A(n1486), .B(n1485), .Y(n442) );
  CLKINVX6TS U530 ( .A(n488), .Y(n487) );
  XOR2X1TS U531 ( .A(n746), .B(n745), .Y(addWeight_26__add_s[3]) );
  NAND2X2TS U532 ( .A(sumOut[97]), .B(n1463), .Y(n1598) );
  NAND2BX2TS U533 ( .AN(sumOut[219]), .B(n623), .Y(n624) );
  NAND2X2TS U534 ( .A(sumOut[208]), .B(n2161), .Y(n740) );
  AOI21X1TS U535 ( .A0(n2267), .A1(n2264), .B0(n2263), .Y(n627) );
  NAND2X4TS U536 ( .A(n657), .B(n1608), .Y(n658) );
  OAI2BB1X2TS U537 ( .A0N(n1502), .A1N(n2005), .B0(n1501), .Y(n1505) );
  NAND2X2TS U538 ( .A(n716), .B(n1666), .Y(n2257) );
  OR2X4TS U539 ( .A(n2380), .B(n725), .Y(n665) );
  OAI21X2TS U540 ( .A0(n1891), .A1(n519), .B0(n1890), .Y(n2222) );
  OAI21X2TS U541 ( .A0(n1836), .A1(n531), .B0(n1835), .Y(n2187) );
  OAI21X2TS U542 ( .A0(n1854), .A1(n487), .B0(n1853), .Y(n2252) );
  BUFX8TS U543 ( .A(n721), .Y(n1670) );
  OAI21X2TS U544 ( .A0(sumOut[3]), .A1(n1519), .B0(n1522), .Y(n476) );
  OAI2BB1X4TS U545 ( .A0N(n1321), .A1N(n1730), .B0(n1320), .Y(n1325) );
  NAND2X2TS U546 ( .A(n2158), .B(n1611), .Y(n587) );
  XOR2X1TS U547 ( .A(n647), .B(n646), .Y(addWeight_27__add_s[6]) );
  OAI2BB1X2TS U548 ( .A0N(n643), .A1N(n599), .B0(n642), .Y(n647) );
  AOI21X2TS U549 ( .A0(n1647), .A1(n1644), .B0(n1643), .Y(n542) );
  OAI2BB1X4TS U550 ( .A0N(n1550), .A1N(n1551), .B0(n1549), .Y(n1555) );
  OAI21X4TS U551 ( .A0(n664), .A1(sumOut[203]), .B0(n665), .Y(n671) );
  XOR2X4TS U552 ( .A(n547), .B(n322), .Y(addWeight_25__add_s[7]) );
  NOR2BX2TS U553 ( .AN(n1566), .B(n546), .Y(n549) );
  CLKAND2X4TS U554 ( .A(sumOut[204]), .B(n1536), .Y(n2015) );
  NOR2X2TS U555 ( .A(n1532), .B(n1533), .Y(n673) );
  AOI21X4TS U556 ( .A0(n2233), .A1(n727), .B0(n726), .Y(n669) );
  NAND2X6TS U557 ( .A(n324), .B(n323), .Y(n727) );
  CLKINVX6TS U558 ( .A(sumOut[203]), .Y(n324) );
  NOR2X4TS U559 ( .A(n1509), .B(n1508), .Y(n1510) );
  NAND2X4TS U560 ( .A(n2017), .B(n1566), .Y(n434) );
  NAND2X4TS U561 ( .A(n434), .B(n1565), .Y(n1570) );
  CLKBUFX2TS U562 ( .A(n2382), .Y(sumOut[200]) );
  NAND2X4TS U563 ( .A(sumOut[248]), .B(n556), .Y(n471) );
  NAND2X4TS U564 ( .A(n470), .B(n471), .Y(n1029) );
  XOR2X4TS U565 ( .A(n1278), .B(n1277), .Y(addWeight_31__add_s[6]) );
  NAND2X4TS U566 ( .A(sumOut[208]), .B(n2161), .Y(n1593) );
  NAND2X4TS U567 ( .A(n1443), .B(n1593), .Y(n1445) );
  NAND2BX2TS U568 ( .AN(n326), .B(n1097), .Y(n1102) );
  NAND2X1TS U569 ( .A(n1096), .B(n1095), .Y(n326) );
  NAND2BX2TS U570 ( .AN(n327), .B(n1057), .Y(n1062) );
  NAND2X1TS U571 ( .A(n1056), .B(n1055), .Y(n327) );
  BUFX6TS U572 ( .A(n2419), .Y(sumOut[88]) );
  AND2X4TS U573 ( .A(n2421), .B(weightsIn[52]), .Y(n2208) );
  AND2X4TS U574 ( .A(n2396), .B(weightsIn[97]), .Y(n2283) );
  NAND2X2TS U575 ( .A(sumOut[128]), .B(n896), .Y(n1872) );
  NAND2X4TS U576 ( .A(n2374), .B(n677), .Y(n332) );
  INVX4TS U577 ( .A(n756), .Y(n543) );
  BUFX8TS U578 ( .A(n756), .Y(n467) );
  OR2X8TS U579 ( .A(n2420), .B(n573), .Y(n704) );
  CLKINVX1TS U580 ( .A(n1880), .Y(sumOut[160]) );
  CLKINVX1TS U581 ( .A(n1945), .Y(sumOut[192]) );
  NOR2X2TS U582 ( .A(n2016), .B(n1532), .Y(n1566) );
  NOR2X2TS U583 ( .A(sumOut[205]), .B(n360), .Y(n1532) );
  OAI2BB1X2TS U584 ( .A0N(n563), .A1N(n599), .B0(n562), .Y(n566) );
  CLKBUFX2TS U585 ( .A(n1729), .Y(n335) );
  CLKBUFX2TS U586 ( .A(n1812), .Y(n336) );
  OAI2BB1X2TS U587 ( .A0N(n1104), .A1N(n1729), .B0(n1106), .Y(n867) );
  NAND2BX4TS U588 ( .AN(n2440), .B(n337), .Y(n1980) );
  NAND2BX4TS U589 ( .AN(n2397), .B(n338), .Y(n1858) );
  NAND2BX4TS U590 ( .AN(n2434), .B(n339), .Y(n1840) );
  NAND2BX4TS U591 ( .AN(n2408), .B(n340), .Y(n1895) );
  NAND2BX4TS U592 ( .AN(n2388), .B(n341), .Y(n1971) );
  NAND2BX4TS U593 ( .AN(n2386), .B(n342), .Y(n1961) );
  NAND2BX4TS U594 ( .AN(n2371), .B(n343), .Y(n1941) );
  NAND2BX4TS U595 ( .AN(n2431), .B(n344), .Y(n1849) );
  NAND2BX4TS U596 ( .AN(n2405), .B(n345), .Y(n1999) );
  NAND2BX4TS U597 ( .AN(n2400), .B(n346), .Y(n1913) );
  NAND2BX4TS U598 ( .AN(n2425), .B(n347), .Y(n1922) );
  NAND2BX4TS U599 ( .AN(n2411), .B(n932), .Y(n1904) );
  NAND2BX4TS U600 ( .AN(n2403), .B(n897), .Y(n1876) );
  BUFX4TS U601 ( .A(n2380), .Y(sumOut[202]) );
  OAI2BB1X4TS U602 ( .A0N(n1363), .A1N(n1777), .B0(n1362), .Y(n1367) );
  OAI2BB1X4TS U603 ( .A0N(n1369), .A1N(n1763), .B0(n1368), .Y(n1373) );
  OAI2BB1X4TS U604 ( .A0N(n1327), .A1N(n1782), .B0(n1326), .Y(n1331) );
  OAI2BB1X4TS U605 ( .A0N(n1309), .A1N(n1721), .B0(n1308), .Y(n1313) );
  OAI2BB1X4TS U606 ( .A0N(n1297), .A1N(n1795), .B0(n1296), .Y(n1301) );
  OAI2BB1X4TS U607 ( .A0N(n1351), .A1N(n1735), .B0(n1350), .Y(n1355) );
  OAI2BB1X4TS U608 ( .A0N(n1315), .A1N(n1748), .B0(n1314), .Y(n1319) );
  OAI2BB1X4TS U609 ( .A0N(n1393), .A1N(n1807), .B0(n1392), .Y(n1397) );
  OAI2BB1X4TS U610 ( .A0N(n1399), .A1N(n1803), .B0(n1398), .Y(n1403) );
  NAND2BX4TS U611 ( .AN(n2428), .B(n969), .Y(n1931) );
  OAI2BB1X4TS U612 ( .A0N(n1339), .A1N(n1772), .B0(n1338), .Y(n1343) );
  OAI2BB1X4TS U613 ( .A0N(n1357), .A1N(n1758), .B0(n1356), .Y(n1361) );
  NAND2BX4TS U614 ( .AN(n2422), .B(n945), .Y(n1831) );
  NAND2BX4TS U615 ( .AN(n2383), .B(n799), .Y(n1951) );
  BUFX4TS U616 ( .A(n2375), .Y(sumOut[233]) );
  AND2X6TS U617 ( .A(n1055), .B(n1053), .Y(n805) );
  NAND2BX4TS U618 ( .AN(n2392), .B(n849), .Y(n1886) );
  NAND2BX4TS U619 ( .AN(n2437), .B(n1006), .Y(n1867) );
  NAND2BX2TS U620 ( .AN(sumOut[94]), .B(n1427), .Y(n1486) );
  OAI2BB1X2TS U621 ( .A0N(n1084), .A1N(n1747), .B0(n1086), .Y(n843) );
  OAI2BB1X2TS U622 ( .A0N(n1387), .A1N(n1747), .B0(n1386), .Y(n1391) );
  OAI2BB1X4TS U623 ( .A0N(n1333), .A1N(n1768), .B0(n1332), .Y(n1337) );
  CLKBUFX2TS U624 ( .A(n1807), .Y(n350) );
  CLKBUFX2TS U625 ( .A(n1803), .Y(n351) );
  CLKBUFX2TS U626 ( .A(n1790), .Y(n352) );
  OAI2BB1X4TS U627 ( .A0N(n1405), .A1N(n1794), .B0(n1404), .Y(n1409) );
  OAI2BB1X2TS U628 ( .A0N(n1234), .A1N(n1795), .B0(n1236), .Y(n1025) );
  OAI2BB1X2TS U629 ( .A0N(n1114), .A1N(n1763), .B0(n1116), .Y(n879) );
  OAI2BB1X2TS U630 ( .A0N(n1214), .A1N(n1721), .B0(n1216), .Y(n1000) );
  OAI2BB1X2TS U631 ( .A0N(n1204), .A1N(n1748), .B0(n1206), .Y(n988) );
  OAI2BB1X2TS U632 ( .A0N(n1144), .A1N(n1735), .B0(n1146), .Y(n915) );
  OAI2BB1X2TS U633 ( .A0N(n1124), .A1N(n1777), .B0(n1126), .Y(n892) );
  OAI2BB1X2TS U634 ( .A0N(n1184), .A1N(n1782), .B0(n1186), .Y(n964) );
  OAI2BB1X2TS U635 ( .A0N(n1164), .A1N(n1772), .B0(n1166), .Y(n939) );
  OAI2BB1X2TS U636 ( .A0N(n1134), .A1N(n1758), .B0(n1136), .Y(n903) );
  OAI2BB1X2TS U637 ( .A0N(n1194), .A1N(n1730), .B0(n1196), .Y(n976) );
  XNOR2X4TS U638 ( .A(n1283), .B(n354), .Y(addWeight_10__add_s[6]) );
  NAND2X2TS U639 ( .A(n1282), .B(n1281), .Y(n354) );
  OAI2BB1X2TS U640 ( .A0N(n1074), .A1N(n1807), .B0(n1076), .Y(n832) );
  OAI2BB1X2TS U641 ( .A0N(n1064), .A1N(n1803), .B0(n1066), .Y(n819) );
  OAI2BB1X2TS U642 ( .A0N(n1044), .A1N(n1790), .B0(n1046), .Y(n793) );
  OAI2BB1X2TS U643 ( .A0N(n1174), .A1N(n1768), .B0(n1176), .Y(n952) );
  OAI2BB1X2TS U644 ( .A0N(n1054), .A1N(n1794), .B0(n1056), .Y(n806) );
  CLKBUFX2TS U645 ( .A(n1811), .Y(n355) );
  NAND2BX2TS U646 ( .AN(n479), .B(n2026), .Y(n478) );
  BUFX4TS U647 ( .A(n2415), .Y(sumOut[97]) );
  OAI2BB1X2TS U648 ( .A0N(n1254), .A1N(n1812), .B0(n1256), .Y(n1252) );
  OAI2BB1X2TS U649 ( .A0N(n697), .A1N(n1812), .B0(n696), .Y(n699) );
  XNOR2X4TS U650 ( .A(n1500), .B(n357), .Y(addWeight_26__add_s[6]) );
  CLKINVX1TS U651 ( .A(n1534), .Y(n358) );
  INVX2TS U652 ( .A(n358), .Y(n359) );
  NAND2BX2TS U653 ( .AN(sumOut[206]), .B(n359), .Y(n1567) );
  CLKINVX1TS U654 ( .A(n1534), .Y(n360) );
  INVX2TS U655 ( .A(weightsIn[1]), .Y(n361) );
  INVX2TS U656 ( .A(weightsIn[11]), .Y(n363) );
  CLKINVX1TS U657 ( .A(weightsIn[135]), .Y(n365) );
  CLKINVX1TS U658 ( .A(n365), .Y(n366) );
  CLKINVX1TS U659 ( .A(n365), .Y(n367) );
  CLKINVX1TS U660 ( .A(weightsIn[81]), .Y(n368) );
  CLKINVX1TS U661 ( .A(n368), .Y(n369) );
  CLKINVX1TS U662 ( .A(n368), .Y(n370) );
  INVX2TS U663 ( .A(weightsIn[16]), .Y(n371) );
  INVX2TS U664 ( .A(weightsIn[76]), .Y(n373) );
  CLKINVX1TS U665 ( .A(n375), .Y(n376) );
  INVX2TS U666 ( .A(n375), .Y(n377) );
  CLKINVX1TS U667 ( .A(n375), .Y(n378) );
  CLKINVX1TS U668 ( .A(n379), .Y(n380) );
  INVX2TS U669 ( .A(n379), .Y(n381) );
  CLKINVX1TS U670 ( .A(n379), .Y(n382) );
  CLKINVX3TS U671 ( .A(weightsIn[98]), .Y(n383) );
  CLKINVX1TS U672 ( .A(n383), .Y(n384) );
  INVX2TS U673 ( .A(n383), .Y(n385) );
  CLKINVX1TS U674 ( .A(n383), .Y(n386) );
  CLKINVX1TS U675 ( .A(n387), .Y(n388) );
  INVX2TS U676 ( .A(n387), .Y(n389) );
  CLKINVX1TS U677 ( .A(n387), .Y(n390) );
  CLKINVX1TS U678 ( .A(n391), .Y(n392) );
  INVX2TS U679 ( .A(n391), .Y(n393) );
  CLKINVX1TS U680 ( .A(n391), .Y(n394) );
  CLKINVX1TS U681 ( .A(weightsIn[136]), .Y(n395) );
  CLKINVX1TS U682 ( .A(n395), .Y(n396) );
  CLKINVX1TS U683 ( .A(n395), .Y(n397) );
  INVX2TS U684 ( .A(weightsIn[21]), .Y(n398) );
  CLKINVX6TS U685 ( .A(n398), .Y(n399) );
  INVX2TS U686 ( .A(weightsIn[26]), .Y(n400) );
  CLKINVX1TS U687 ( .A(n400), .Y(n401) );
  INVX2TS U688 ( .A(weightsIn[31]), .Y(n403) );
  CLKINVX6TS U689 ( .A(n403), .Y(n404) );
  INVX2TS U690 ( .A(weightsIn[36]), .Y(n405) );
  CLKINVX6TS U691 ( .A(n405), .Y(n406) );
  INVX2TS U692 ( .A(weightsIn[41]), .Y(n407) );
  CLKINVX6TS U693 ( .A(n407), .Y(n408) );
  INVX2TS U694 ( .A(weightsIn[46]), .Y(n409) );
  CLKINVX6TS U695 ( .A(n409), .Y(n410) );
  INVX2TS U696 ( .A(weightsIn[66]), .Y(n411) );
  CLKINVX6TS U697 ( .A(n411), .Y(n412) );
  INVX2TS U698 ( .A(weightsIn[71]), .Y(n413) );
  INVX2TS U699 ( .A(weightsIn[86]), .Y(n415) );
  CLKINVX6TS U700 ( .A(n415), .Y(n416) );
  INVX2TS U701 ( .A(weightsIn[91]), .Y(n417) );
  CLKINVX1TS U702 ( .A(n417), .Y(n418) );
  NAND2X2TS U703 ( .A(n2404), .B(n369), .Y(n491) );
  INVX2TS U704 ( .A(n1573), .Y(n480) );
  NAND2X1TS U705 ( .A(n643), .B(n644), .Y(n600) );
  INVX2TS U706 ( .A(n742), .Y(n1440) );
  OR2X4TS U707 ( .A(n2441), .B(n372), .Y(n536) );
  OR2X4TS U708 ( .A(n2406), .B(n374), .Y(n518) );
  CLKBUFX2TS U709 ( .A(weightsIn[131]), .Y(n1442) );
  CLKBUFX2TS U710 ( .A(weightsIn[61]), .Y(n1463) );
  CLKBUFX2TS U711 ( .A(weightsIn[146]), .Y(n733) );
  NAND2X1TS U712 ( .A(n1279), .B(n1282), .Y(n580) );
  NOR2X1TS U713 ( .A(sumOut[141]), .B(n1130), .Y(n1365) );
  INVX2TS U714 ( .A(sumOut[80]), .Y(n700) );
  OR2X4TS U715 ( .A(n2448), .B(n362), .Y(n1521) );
  INVX2TS U716 ( .A(n1607), .Y(n773) );
  NOR2X1TS U717 ( .A(n1538), .B(n1544), .Y(n1491) );
  OAI2BB1X2TS U718 ( .A0N(n1479), .A1N(n1560), .B0(n1478), .Y(n1483) );
  OAI2BB1X2TS U719 ( .A0N(n1224), .A1N(n1717), .B0(n1226), .Y(n1013) );
  OAI2BB1X2TS U720 ( .A0N(n1154), .A1N(n1753), .B0(n1156), .Y(n927) );
  OAI2BB1X2TS U721 ( .A0N(n1264), .A1N(n1811), .B0(n1266), .Y(n1247) );
  AOI21X1TS U722 ( .A0(n2252), .A1(n2249), .B0(n2248), .Y(n1861) );
  AOI21X1TS U723 ( .A0(n2222), .A1(n2219), .B0(n2218), .Y(n1898) );
  AOI21X1TS U724 ( .A0(n2187), .A1(n2184), .B0(n2183), .Y(n1843) );
  AOI21X1TS U725 ( .A0(n2282), .A1(n2279), .B0(n2278), .Y(n1993) );
  OAI2BB1X2TS U726 ( .A0N(n1094), .A1N(n1743), .B0(n1096), .Y(n856) );
  XOR2X1TS U727 ( .A(n780), .B(n779), .Y(addWeight_1__add_s[3]) );
  OR2X4TS U728 ( .A(sumOut[17]), .B(n364), .Y(n1611) );
  OAI2BB1X2TS U729 ( .A0N(n1507), .A1N(n2005), .B0(n1506), .Y(n1511) );
  NAND2X2TS U730 ( .A(n478), .B(n477), .Y(n1531) );
  AND2X4TS U731 ( .A(n1571), .B(n1574), .Y(n477) );
  NOR2X2TS U732 ( .A(n1544), .B(n1543), .Y(n1545) );
  INVX1TS U733 ( .A(n2016), .Y(n672) );
  NAND2X2TS U734 ( .A(n481), .B(n1527), .Y(n1573) );
  NOR2X4TS U735 ( .A(n1514), .B(n2007), .Y(n1496) );
  NAND2X2TS U736 ( .A(sumOut[169]), .B(n1663), .Y(n1986) );
  NAND2X2TS U737 ( .A(sumOut[177]), .B(n1691), .Y(n1967) );
  NAND2X2TS U738 ( .A(sumOut[185]), .B(n1704), .Y(n1957) );
  NAND2X2TS U739 ( .A(sumOut[193]), .B(n1654), .Y(n1947) );
  NAND2X2TS U740 ( .A(sumOut[241]), .B(n1709), .Y(n1937) );
  INVX3TS U741 ( .A(n1599), .Y(n747) );
  NAND2X2TS U742 ( .A(sumOut[249]), .B(n555), .Y(n1666) );
  NAND2X2TS U743 ( .A(sumOut[161]), .B(n1673), .Y(n1882) );
  AND2X4TS U744 ( .A(sumOut[148]), .B(n1120), .Y(n1764) );
  AND2X4TS U745 ( .A(sumOut[44]), .B(n1220), .Y(n1722) );
  AND2X4TS U746 ( .A(sumOut[140]), .B(n1130), .Y(n1778) );
  AND2X4TS U747 ( .A(sumOut[60]), .B(n1200), .Y(n1731) );
  AND2X4TS U748 ( .A(sumOut[76]), .B(n1180), .Y(n1769) );
  AND2X4TS U749 ( .A(sumOut[108]), .B(n1170), .Y(n1773) );
  AND2X4TS U750 ( .A(sumOut[52]), .B(n1210), .Y(n1749) );
  AND2X4TS U751 ( .A(sumOut[28]), .B(n1240), .Y(n1796) );
  AND2X4TS U752 ( .A(sumOut[124]), .B(n1150), .Y(n1736) );
  AND2X4TS U753 ( .A(sumOut[132]), .B(n1140), .Y(n1759) );
  AND2X4TS U754 ( .A(sumOut[68]), .B(n1190), .Y(n1783) );
  AND2X4TS U755 ( .A(sumOut[36]), .B(n1230), .Y(n1718) );
  AND2X4TS U756 ( .A(sumOut[116]), .B(n1160), .Y(n1754) );
  AND2X4TS U757 ( .A(sumOut[188]), .B(n1070), .Y(n1800) );
  AND2X4TS U758 ( .A(sumOut[180]), .B(n1080), .Y(n1804) );
  AND2X4TS U759 ( .A(sumOut[20]), .B(n1260), .Y(n1813) );
  INVX2TS U760 ( .A(n751), .Y(n468) );
  AND2X4TS U761 ( .A(sumOut[172]), .B(n1090), .Y(n1744) );
  INVX2TS U762 ( .A(n743), .Y(n473) );
  AND2X4TS U763 ( .A(sumOut[244]), .B(n1050), .Y(n1787) );
  AND2X4TS U764 ( .A(sumOut[196]), .B(n1060), .Y(n1791) );
  AND2X4TS U765 ( .A(sumOut[164]), .B(n1100), .Y(n1740) );
  NAND2X2TS U766 ( .A(sumOut[221]), .B(n603), .Y(n601) );
  AND2X4TS U767 ( .A(sumOut[228]), .B(n1437), .Y(n1557) );
  INVX2TS U768 ( .A(n1026), .Y(n463) );
  INVX3TS U769 ( .A(sumOut[6]), .Y(n481) );
  INVX4TS U770 ( .A(n872), .Y(n873) );
  INVX2TS U771 ( .A(n577), .Y(n579) );
  INVX4TS U772 ( .A(n920), .Y(n921) );
  INVX4TS U773 ( .A(n825), .Y(n826) );
  INVX4TS U774 ( .A(n812), .Y(n813) );
  INVX2TS U775 ( .A(n857), .Y(n865) );
  INVX4TS U776 ( .A(n885), .Y(n886) );
  INVX4TS U777 ( .A(n908), .Y(n909) );
  INVX4TS U778 ( .A(n993), .Y(n994) );
  INVX4TS U779 ( .A(n1018), .Y(n1019) );
  INVX4TS U780 ( .A(n786), .Y(n787) );
  INVX4TS U781 ( .A(n957), .Y(n958) );
  INVX4TS U782 ( .A(n981), .Y(n982) );
  BUFX4TS U783 ( .A(weightsIn[147]), .Y(n677) );
  NAND2BX2TS U784 ( .AN(n464), .B(n1453), .Y(n1458) );
  XOR2X1TS U785 ( .A(n754), .B(n753), .Y(addWeight_12__add_s[3]) );
  AOI21X2TS U786 ( .A0(n1632), .A1(n1629), .B0(n1628), .Y(n746) );
  XOR2X2TS U787 ( .A(n771), .B(n770), .Y(addWeight_11__add_s[3]) );
  AOI21X1TS U788 ( .A0(n2247), .A1(n2244), .B0(n2243), .Y(n1889) );
  AOI21X1TS U789 ( .A0(n2277), .A1(n2274), .B0(n2273), .Y(n1964) );
  AOI21X1TS U790 ( .A0(n2242), .A1(n2239), .B0(n2238), .Y(n1954) );
  AOI21X1TS U791 ( .A0(n2262), .A1(n2259), .B0(n2258), .Y(n1944) );
  NAND2X4TS U792 ( .A(n587), .B(n1610), .Y(n2297) );
  AOI21X1TS U793 ( .A0(n2292), .A1(n2289), .B0(n2288), .Y(n1974) );
  NAND2X4TS U794 ( .A(n492), .B(n516), .Y(n445) );
  NAND2X2TS U795 ( .A(n741), .B(n1592), .Y(n1632) );
  AOI2BB1X2TS U796 ( .A0N(sumOut[56]), .A1N(n968), .B0(n635), .Y(
        addWeight_7__add_s[0]) );
  AOI2BB1X2TS U797 ( .A0N(sumOut[120]), .A1N(n907), .B0(n636), .Y(
        addWeight_15__add_s[0]) );
  AOI2BB1X2TS U798 ( .A0N(sumOut[72]), .A1N(n943), .B0(n637), .Y(
        addWeight_9__add_s[0]) );
  AOI2BB1X2TS U799 ( .A0N(sumOut[48]), .A1N(n980), .B0(n638), .Y(
        addWeight_6__add_s[0]) );
  AOI2BB1X2TS U800 ( .A0N(sumOut[64]), .A1N(n956), .B0(n639), .Y(
        addWeight_8__add_s[0]) );
  AOI2BB1X2TS U801 ( .A0N(sumOut[136]), .A1N(n883), .B0(n640), .Y(
        addWeight_17__add_s[0]) );
  AOI2BB1X2TS U802 ( .A0N(sumOut[104]), .A1N(n931), .B0(n634), .Y(
        addWeight_13__add_s[0]) );
  AOI2BB1X2TS U803 ( .A0N(sumOut[8]), .A1N(n2170), .B0(n2169), .Y(
        addWeight_1__add_s[0]) );
  AOI2BB1X2TS U804 ( .A0N(sumOut[88]), .A1N(n2167), .B0(n2166), .Y(
        addWeight_11__add_s[0]) );
  AOI2BB1X2TS U805 ( .A0N(sumOut[112]), .A1N(n919), .B0(n633), .Y(
        addWeight_14__add_s[0]) );
  AOI2BB1X2TS U806 ( .A0N(sumOut[32]), .A1N(n1004), .B0(n631), .Y(
        addWeight_4__add_s[0]) );
  AOI2BB1X2TS U807 ( .A0N(sumOut[144]), .A1N(n871), .B0(n632), .Y(
        addWeight_18__add_s[0]) );
  AOI2BB1X2TS U808 ( .A0N(sumOut[40]), .A1N(n992), .B0(n630), .Y(
        addWeight_5__add_s[0]) );
  AOI2BB1X2TS U809 ( .A0N(sumOut[24]), .A1N(n1017), .B0(n629), .Y(
        addWeight_3__add_s[0]) );
  NAND2X4TS U810 ( .A(n1700), .B(n491), .Y(n492) );
  NAND2X4TS U811 ( .A(n1702), .B(n484), .Y(n486) );
  NAND2X4TS U812 ( .A(n1657), .B(n482), .Y(n483) );
  NAND2X4TS U813 ( .A(n1685), .B(n504), .Y(n505) );
  NAND2X4TS U814 ( .A(n1689), .B(n506), .Y(n507) );
  NAND2X2TS U815 ( .A(n1504), .B(n1503), .Y(n551) );
  NAND2X4TS U816 ( .A(n1687), .B(n510), .Y(n512) );
  NAND2X4TS U817 ( .A(n1678), .B(n513), .Y(n514) );
  NAND2X4TS U818 ( .A(n1698), .B(n508), .Y(n509) );
  NAND2X4TS U819 ( .A(n1676), .B(n499), .Y(n501) );
  NAND2X4TS U820 ( .A(n1715), .B(n502), .Y(n503) );
  NAND2X4TS U821 ( .A(n1707), .B(n493), .Y(n494) );
  NAND2X4TS U822 ( .A(n1680), .B(n495), .Y(n496) );
  NAND2X4TS U823 ( .A(n1652), .B(n497), .Y(n498) );
  NAND2X2TS U824 ( .A(n1956), .B(n2143), .Y(n1958) );
  NAND2X2TS U825 ( .A(n1966), .B(n2147), .Y(n1968) );
  NAND2X2TS U826 ( .A(n1985), .B(n2149), .Y(n1987) );
  NAND2X2TS U827 ( .A(n1881), .B(n2154), .Y(n1883) );
  NAND2X2TS U828 ( .A(n1936), .B(n2156), .Y(n1938) );
  NAND2X2TS U829 ( .A(n1946), .B(n2137), .Y(n1948) );
  NAND2X2TS U830 ( .A(n1817), .B(n2139), .Y(n1819) );
  OAI21X2TS U831 ( .A0(n748), .A1(n747), .B0(n1598), .Y(n1642) );
  NAND2X2TS U832 ( .A(n715), .B(n1667), .Y(n716) );
  NAND2BX2TS U833 ( .AN(n527), .B(n1926), .Y(n1686) );
  NAND2BX2TS U834 ( .AN(n521), .B(n1899), .Y(n1653) );
  NAND2BX2TS U835 ( .AN(n517), .B(n1994), .Y(n1708) );
  NAND2BX2TS U836 ( .AN(n519), .B(n1890), .Y(n1681) );
  NAND2BX2TS U837 ( .AN(n487), .B(n1853), .Y(n1658) );
  NAND2BX2TS U838 ( .AN(n533), .B(n1862), .Y(n1688) );
  NAND2BX2TS U839 ( .AN(n523), .B(n1826), .Y(n1677) );
  NAND2BX2TS U840 ( .AN(n531), .B(n1835), .Y(n1699) );
  NAND2BX2TS U841 ( .AN(n529), .B(n1844), .Y(n1690) );
  NAND2BX2TS U842 ( .AN(n535), .B(n1975), .Y(n1679) );
  NAND2BX2TS U843 ( .AN(n515), .B(n1871), .Y(n1701) );
  NAND2BX2TS U844 ( .AN(n525), .B(n1917), .Y(n1716) );
  NAND2BX2TS U845 ( .AN(n489), .B(n1908), .Y(n1703) );
  NAND2X4TS U846 ( .A(n931), .B(n2413), .Y(n1652) );
  NAND2X4TS U847 ( .A(n956), .B(n2427), .Y(n1715) );
  NAND2X4TS U848 ( .A(n907), .B(n2407), .Y(n1707) );
  NOR2X2TS U849 ( .A(n1346), .B(n1754), .Y(n1156) );
  NOR2X2TS U850 ( .A(n1352), .B(n1736), .Y(n1146) );
  NAND2X4TS U851 ( .A(n485), .B(n2402), .Y(n1702) );
  NOR2X2TS U852 ( .A(n1334), .B(n1769), .Y(n1176) );
  NAND2X4TS U853 ( .A(n500), .B(n2424), .Y(n1676) );
  NAND2X4TS U854 ( .A(n919), .B(n2410), .Y(n1680) );
  NAND2X4TS U855 ( .A(n896), .B(sumOut[128]), .Y(n1700) );
  NOR2X2TS U856 ( .A(n1298), .B(n1796), .Y(n1236) );
  NAND2X4TS U857 ( .A(n1017), .B(n2442), .Y(n1678) );
  NOR2X2TS U858 ( .A(n1406), .B(n1791), .Y(n1056) );
  NOR2X2TS U859 ( .A(n1304), .B(n1718), .Y(n1226) );
  NAND2X4TS U860 ( .A(n511), .B(n2439), .Y(n1687) );
  NOR2X2TS U861 ( .A(n1310), .B(n1722), .Y(n1216) );
  NAND2X4TS U862 ( .A(n992), .B(n2436), .Y(n1698) );
  NOR2X2TS U863 ( .A(n1382), .B(n1740), .Y(n1096) );
  NAND2X4TS U864 ( .A(n980), .B(n2433), .Y(n1689) );
  NAND2X4TS U865 ( .A(n968), .B(n2430), .Y(n1685) );
  NAND2X4TS U866 ( .A(n871), .B(n2399), .Y(n1657) );
  INVX1TS U867 ( .A(n1556), .Y(n1559) );
  INVX1TS U868 ( .A(n1538), .Y(n1541) );
  INVX1TS U869 ( .A(n1547), .Y(n1550) );
  INVX1TS U870 ( .A(n617), .Y(n563) );
  INVX1TS U871 ( .A(n1809), .Y(n683) );
  NOR2X2TS U872 ( .A(n1287), .B(n1286), .Y(n1288) );
  INVX1TS U873 ( .A(n2011), .Y(n1285) );
  INVX2TS U874 ( .A(n2023), .Y(n1578) );
  NOR2X2TS U875 ( .A(n1508), .B(n2003), .Y(n1501) );
  INVX1TS U876 ( .A(n2019), .Y(n1291) );
  NAND2X2TS U877 ( .A(sumOut[89]), .B(n763), .Y(n1602) );
  NAND2X2TS U878 ( .A(sumOut[9]), .B(n772), .Y(n1606) );
  INVX2TS U879 ( .A(n608), .Y(n715) );
  CLKINVX2TS U880 ( .A(n1567), .Y(n546) );
  NAND2X4TS U881 ( .A(n537), .B(n538), .Y(n777) );
  NAND2X4TS U882 ( .A(n539), .B(n540), .Y(n768) );
  NAND2X2TS U883 ( .A(sumOut[201]), .B(n723), .Y(n1669) );
  NAND2X2TS U884 ( .A(n1520), .B(n1713), .Y(n1522) );
  NOR2X1TS U885 ( .A(sumOut[223]), .B(n603), .Y(n604) );
  AND2X2TS U886 ( .A(sumOut[229]), .B(n1433), .Y(n1561) );
  AND2X4TS U887 ( .A(sumOut[220]), .B(n605), .Y(n618) );
  AND2X4TS U888 ( .A(sumOut[84]), .B(n584), .Y(n2020) );
  INVX2TS U889 ( .A(n1451), .Y(n1452) );
  INVX2TS U890 ( .A(n1470), .Y(n1471) );
  INVX2TS U891 ( .A(n682), .Y(n1245) );
  CLKINVX2TS U892 ( .A(n1432), .Y(n1433) );
  INVX2TS U893 ( .A(n893), .Y(n901) );
  INVX2TS U894 ( .A(n880), .Y(n890) );
  INVX3TS U895 ( .A(n883), .Y(n884) );
  INVX2TS U896 ( .A(n868), .Y(n877) );
  INVX2TS U897 ( .A(n844), .Y(n854) );
  INVX2TS U898 ( .A(n953), .Y(n962) );
  INVX2TS U899 ( .A(n940), .Y(n950) );
  INVX3TS U900 ( .A(n943), .Y(n944) );
  INVX2TS U901 ( .A(n928), .Y(n937) );
  INVX2TS U902 ( .A(n1461), .Y(n1462) );
  INVX2TS U903 ( .A(n916), .Y(n925) );
  INVX2TS U904 ( .A(n904), .Y(n913) );
  INVX2TS U905 ( .A(n1424), .Y(n1425) );
  INVX2TS U906 ( .A(n1416), .Y(n1417) );
  INVX2TS U907 ( .A(n695), .Y(n1250) );
  INVX2TS U908 ( .A(n833), .Y(n841) );
  INVX2TS U909 ( .A(n820), .Y(n830) );
  INVX2TS U910 ( .A(n807), .Y(n817) );
  INVX2TS U911 ( .A(n794), .Y(n804) );
  INVX2TS U912 ( .A(n781), .Y(n791) );
  INVX2TS U913 ( .A(n989), .Y(n998) );
  INVX2TS U914 ( .A(n1014), .Y(n1023) );
  INVX2TS U915 ( .A(n977), .Y(n986) );
  INVX3TS U916 ( .A(n1004), .Y(n1005) );
  INVX2TS U917 ( .A(n965), .Y(n974) );
  INVX2TS U918 ( .A(n1001), .Y(n1011) );
  BUFX3TS U919 ( .A(weightsIn[116]), .Y(n1704) );
  BUFX3TS U920 ( .A(weightsIn[56]), .Y(n763) );
  BUFX4TS U921 ( .A(weightsIn[32]), .Y(n978) );
  BUFX4TS U922 ( .A(weightsIn[67]), .Y(n929) );
  BUFX3TS U923 ( .A(weightsIn[151]), .Y(n1709) );
  BUFX3TS U924 ( .A(weightsIn[126]), .Y(n723) );
  BUFX3TS U925 ( .A(weightsIn[121]), .Y(n1654) );
  BUFX3TS U926 ( .A(weightsIn[10]), .Y(n2159) );
  BUFX4TS U927 ( .A(weightsIn[42]), .Y(n954) );
  BUFX4TS U928 ( .A(weightsIn[37]), .Y(n966) );
  BUFX3TS U929 ( .A(weightsIn[130]), .Y(n2161) );
  BUFX3TS U930 ( .A(weightsIn[6]), .Y(n772) );
  BUFX4TS U931 ( .A(weightsIn[47]), .Y(n941) );
  BUFX4TS U932 ( .A(weightsIn[22]), .Y(n1002) );
  BUFX3TS U933 ( .A(weightsIn[141]), .Y(n755) );
  BUFX3TS U934 ( .A(weightsIn[106]), .Y(n1663) );
  BUFX4TS U935 ( .A(weightsIn[87]), .Y(n881) );
  BUFX3TS U936 ( .A(weightsIn[101]), .Y(n1673) );
  BUFX4TS U937 ( .A(weightsIn[82]), .Y(n894) );
  BUFX3TS U938 ( .A(weightsIn[111]), .Y(n1691) );
  INVX2TS U939 ( .A(weightsIn[12]), .Y(n420) );
  OAI21X4TS U940 ( .A0(n1033), .A1(n1034), .B0(n1032), .Y(n2014) );
  BUFX4TS U941 ( .A(n2370), .Y(sumOut[249]) );
  BUFX6TS U942 ( .A(n2442), .Y(sumOut[24]) );
  BUFX6TS U943 ( .A(n2436), .Y(sumOut[40]) );
  BUFX6TS U944 ( .A(n2439), .Y(sumOut[32]) );
  BUFX6TS U945 ( .A(n2399), .Y(sumOut[144]) );
  BUFX6TS U946 ( .A(n2410), .Y(sumOut[112]) );
  BUFX6TS U947 ( .A(n2413), .Y(sumOut[104]) );
  BUFX6TS U948 ( .A(n2430), .Y(sumOut[56]) );
  BUFX6TS U949 ( .A(n2407), .Y(sumOut[120]) );
  BUFX6TS U950 ( .A(n2424), .Y(sumOut[72]) );
  BUFX6TS U951 ( .A(n2433), .Y(sumOut[48]) );
  BUFX6TS U952 ( .A(n2427), .Y(sumOut[64]) );
  BUFX6TS U953 ( .A(n2402), .Y(sumOut[136]) );
  NAND2BX4TS U954 ( .AN(sumOut[18]), .B(n420), .Y(n687) );
  OAI21X4TS U955 ( .A0(n670), .A1(n671), .B0(n669), .Y(n2017) );
  BUFX3TS U956 ( .A(n2381), .Y(sumOut[201]) );
  BUFX3TS U957 ( .A(n2391), .Y(sumOut[169]) );
  BUFX3TS U958 ( .A(n2389), .Y(sumOut[177]) );
  BUFX3TS U959 ( .A(n2384), .Y(sumOut[193]) );
  BUFX3TS U960 ( .A(n2387), .Y(sumOut[185]) );
  BUFX3TS U961 ( .A(n2372), .Y(sumOut[241]) );
  BUFX3TS U962 ( .A(n2393), .Y(sumOut[161]) );
  NAND2X2TS U963 ( .A(n1551), .B(n442), .Y(n1426) );
  BUFX3TS U964 ( .A(n2445), .Y(sumOut[9]) );
  BUFX3TS U965 ( .A(n2418), .Y(sumOut[89]) );
  OAI21X4TS U966 ( .A0(n900), .A1(n445), .B0(n899), .Y(n1758) );
  NAND2X2TS U967 ( .A(n447), .B(n1577), .Y(n1582) );
  NAND2X2TS U968 ( .A(n2026), .B(n1578), .Y(n447) );
  BUFX3TS U969 ( .A(n2448), .Y(sumOut[1]) );
  BUFX6TS U970 ( .A(n2435), .Y(sumOut[41]) );
  BUFX6TS U971 ( .A(n2438), .Y(sumOut[33]) );
  BUFX6TS U972 ( .A(n2398), .Y(sumOut[145]) );
  BUFX6TS U973 ( .A(n2409), .Y(sumOut[113]) );
  BUFX6TS U974 ( .A(n2412), .Y(sumOut[105]) );
  BUFX6TS U975 ( .A(n2429), .Y(sumOut[57]) );
  BUFX6TS U976 ( .A(n2423), .Y(sumOut[73]) );
  BUFX6TS U977 ( .A(n2432), .Y(sumOut[49]) );
  BUFX6TS U978 ( .A(n2426), .Y(sumOut[65]) );
  BUFX6TS U979 ( .A(n2401), .Y(sumOut[137]) );
  XNOR2X4TS U980 ( .A(n461), .B(n673), .Y(addWeight_25__add_s[5]) );
  AOI21X4TS U981 ( .A0(n2017), .A1(n672), .B0(n2015), .Y(n461) );
  NAND2BX2TS U982 ( .AN(n1454), .B(sumOut[214]), .Y(n1499) );
  BUFX6TS U983 ( .A(n2293), .Y(n462) );
  NAND2BX4TS U984 ( .AN(n2369), .B(n463), .Y(n1031) );
  OAI2BB1X4TS U985 ( .A0N(n688), .A1N(n689), .B0(n1611), .Y(n693) );
  XOR2X4TS U986 ( .A(n1495), .B(n1494), .Y(addWeight_1__add_s[6]) );
  XOR2X4TS U987 ( .A(n1489), .B(n1488), .Y(addWeight_11__add_s[6]) );
  XOR2X4TS U988 ( .A(n1252), .B(n1251), .Y(addWeight_2__add_s[6]) );
  XOR2X4TS U989 ( .A(n699), .B(n698), .Y(addWeight_2__add_s[5]) );
  OR2X8TS U990 ( .A(n2381), .B(n723), .Y(n721) );
  NAND2BX2TS U991 ( .AN(n465), .B(n1418), .Y(n1423) );
  NAND2X1TS U992 ( .A(n1490), .B(n1493), .Y(n465) );
  NAND2X1TS U993 ( .A(n1484), .B(n1487), .Y(n466) );
  NOR2X2TS U994 ( .A(n1244), .B(n1808), .Y(n1266) );
  NAND2BX4TS U995 ( .AN(n2414), .B(n468), .Y(n1466) );
  NAND2X4TS U996 ( .A(n2381), .B(n723), .Y(n666) );
  BUFX6TS U997 ( .A(n2416), .Y(sumOut[96]) );
  NAND2X4TS U998 ( .A(sumOut[225]), .B(n755), .Y(n610) );
  OAI2BB1X4TS U999 ( .A0N(n1695), .A1N(n675), .B0(n731), .Y(n680) );
  XOR2X4TS U1000 ( .A(n867), .B(n866), .Y(addWeight_19__add_s[6]) );
  XOR2X4TS U1001 ( .A(n1483), .B(n1482), .Y(addWeight_28__add_s[6]) );
  OAI2BB1X4TS U1002 ( .A0N(n1682), .A1N(sumOut[153]), .B0(n1683), .Y(n860) );
  NAND2X4TS U1003 ( .A(n860), .B(n1817), .Y(n863) );
  XOR2X4TS U1004 ( .A(n1247), .B(n1246), .Y(addWeight_29__add_s[6]) );
  NAND2X4TS U1005 ( .A(n2370), .B(n555), .Y(n470) );
  NAND2BX4TS U1006 ( .AN(sumOut[210]), .B(n742), .Y(n1441) );
  NAND2X4TS U1007 ( .A(n1661), .B(n472), .Y(n558) );
  NAND2X4TS U1008 ( .A(sumOut[217]), .B(n397), .Y(n472) );
  NAND2X4TS U1009 ( .A(sumOut[216]), .B(n366), .Y(n1661) );
  NAND2BX4TS U1010 ( .AN(n2379), .B(n473), .Y(n1447) );
  OAI21X4TS U1011 ( .A0(n476), .A1(n475), .B0(n474), .Y(n2026) );
  AOI21X4TS U1012 ( .A0(n1618), .A1(n1524), .B0(n1523), .Y(n474) );
  NAND2X4TS U1013 ( .A(n2382), .B(n2146), .Y(n1671) );
  NAND2X4TS U1014 ( .A(n666), .B(n1671), .Y(n667) );
  XOR2X4TS U1015 ( .A(n843), .B(n842), .Y(addWeight_21__add_s[6]) );
  XOR2X4TS U1016 ( .A(n1576), .B(n1575), .Y(addWeight_0__add_s[6]) );
  XOR2X4TS U1017 ( .A(n1025), .B(n1024), .Y(addWeight_3__add_s[6]) );
  XOR2X4TS U1018 ( .A(n1013), .B(n1012), .Y(addWeight_4__add_s[6]) );
  XOR2X4TS U1019 ( .A(n793), .B(n792), .Y(addWeight_30__add_s[6]) );
  XOR2X4TS U1020 ( .A(n806), .B(n805), .Y(addWeight_24__add_s[6]) );
  XOR2X4TS U1021 ( .A(n819), .B(n818), .Y(addWeight_23__add_s[6]) );
  XOR2X4TS U1022 ( .A(n832), .B(n831), .Y(addWeight_22__add_s[6]) );
  XOR2X4TS U1023 ( .A(n856), .B(n855), .Y(addWeight_20__add_s[6]) );
  NAND2X4TS U1024 ( .A(n488), .B(n483), .Y(n875) );
  NAND2X4TS U1025 ( .A(n490), .B(n486), .Y(n888) );
  NAND2X4TS U1026 ( .A(n518), .B(n494), .Y(n911) );
  NAND2X4TS U1027 ( .A(n520), .B(n496), .Y(n923) );
  NAND2X4TS U1028 ( .A(n522), .B(n498), .Y(n935) );
  NAND2X4TS U1029 ( .A(n524), .B(n501), .Y(n948) );
  NAND2X4TS U1030 ( .A(n526), .B(n503), .Y(n960) );
  NAND2X4TS U1031 ( .A(n528), .B(n505), .Y(n972) );
  NAND2X4TS U1032 ( .A(n530), .B(n507), .Y(n984) );
  NAND2X4TS U1033 ( .A(n532), .B(n509), .Y(n996) );
  NAND2X4TS U1034 ( .A(n534), .B(n512), .Y(n1009) );
  NAND2X4TS U1035 ( .A(n536), .B(n514), .Y(n1021) );
  BUFX8TS U1036 ( .A(n2447), .Y(sumOut[3]) );
  XOR2X4TS U1037 ( .A(n1000), .B(n999), .Y(addWeight_5__add_s[6]) );
  XOR2X4TS U1038 ( .A(n988), .B(n987), .Y(addWeight_6__add_s[6]) );
  XOR2X4TS U1039 ( .A(n976), .B(n975), .Y(addWeight_7__add_s[6]) );
  XOR2X4TS U1040 ( .A(n964), .B(n963), .Y(addWeight_8__add_s[6]) );
  XOR2X4TS U1041 ( .A(n952), .B(n951), .Y(addWeight_9__add_s[6]) );
  XOR2X4TS U1042 ( .A(n939), .B(n938), .Y(addWeight_13__add_s[6]) );
  XOR2X4TS U1043 ( .A(n927), .B(n926), .Y(addWeight_14__add_s[6]) );
  XOR2X4TS U1044 ( .A(n915), .B(n914), .Y(addWeight_15__add_s[6]) );
  XOR2X4TS U1045 ( .A(n903), .B(n902), .Y(addWeight_16__add_s[6]) );
  XOR2X4TS U1046 ( .A(n892), .B(n891), .Y(addWeight_17__add_s[6]) );
  XOR2X4TS U1047 ( .A(n879), .B(n878), .Y(addWeight_18__add_s[6]) );
  NAND2X4TS U1048 ( .A(n2398), .B(n419), .Y(n482) );
  OR2X8TS U1049 ( .A(n2398), .B(n418), .Y(n488) );
  NAND2X4TS U1050 ( .A(n2401), .B(n416), .Y(n484) );
  OR2X8TS U1051 ( .A(n2401), .B(n416), .Y(n490) );
  INVX2TS U1052 ( .A(n490), .Y(n489) );
  OR2X8TS U1053 ( .A(n2404), .B(n370), .Y(n516) );
  NAND2X4TS U1054 ( .A(n2409), .B(n414), .Y(n495) );
  NAND2X4TS U1055 ( .A(n2412), .B(n412), .Y(n497) );
  OR2X8TS U1056 ( .A(n2412), .B(n412), .Y(n522) );
  NAND2X4TS U1057 ( .A(n2423), .B(n410), .Y(n499) );
  OR2X8TS U1058 ( .A(n2423), .B(n410), .Y(n524) );
  NAND2X4TS U1059 ( .A(n2426), .B(n408), .Y(n502) );
  OR2X8TS U1060 ( .A(n2426), .B(n408), .Y(n526) );
  NAND2X4TS U1061 ( .A(n2429), .B(n406), .Y(n504) );
  OR2X8TS U1062 ( .A(n2429), .B(n406), .Y(n528) );
  NAND2X4TS U1063 ( .A(n2432), .B(n404), .Y(n506) );
  OR2X8TS U1064 ( .A(n2432), .B(n404), .Y(n530) );
  NAND2X4TS U1065 ( .A(n2435), .B(n402), .Y(n508) );
  NAND2X4TS U1066 ( .A(n2438), .B(n399), .Y(n510) );
  OR2X8TS U1067 ( .A(n2438), .B(n399), .Y(n534) );
  INVX2TS U1068 ( .A(n516), .Y(n515) );
  INVX2TS U1069 ( .A(n522), .Y(n521) );
  INVX2TS U1070 ( .A(n524), .Y(n523) );
  INVX2TS U1071 ( .A(n526), .Y(n525) );
  INVX2TS U1072 ( .A(n528), .Y(n527) );
  INVX2TS U1073 ( .A(n530), .Y(n529) );
  INVX2TS U1074 ( .A(n534), .Y(n533) );
  CLKINVX3TS U1075 ( .A(n2444), .Y(n537) );
  INVX2TS U1076 ( .A(n377), .Y(n538) );
  CLKINVX3TS U1077 ( .A(n2417), .Y(n539) );
  INVX2TS U1078 ( .A(n381), .Y(n540) );
  NAND2BX4TS U1079 ( .AN(n2377), .B(n541), .Y(n760) );
  INVX2TS U1080 ( .A(n393), .Y(n541) );
  NAND2BXLTS U1081 ( .AN(n467), .B(n1595), .Y(n1597) );
  NAND2X4TS U1082 ( .A(n611), .B(n543), .Y(n614) );
  NOR2X4TS U1083 ( .A(sumOut[225]), .B(n755), .Y(n756) );
  NAND2BX4TS U1084 ( .AN(n2390), .B(n544), .Y(n1990) );
  INVX2TS U1085 ( .A(n389), .Y(n544) );
  NAND2BX4TS U1086 ( .AN(n2395), .B(n545), .Y(n1822) );
  INVX2TS U1087 ( .A(n385), .Y(n545) );
  AOI21X4TS U1088 ( .A0(n2017), .A1(n549), .B0(n548), .Y(n547) );
  INVX2TS U1089 ( .A(weightsIn[129]), .Y(n1534) );
  NAND2X4TS U1090 ( .A(n1445), .B(n1444), .Y(n1449) );
  NAND2BX2TS U1091 ( .AN(sumOut[86]), .B(n582), .Y(n1281) );
  OAI21X4TS U1092 ( .A0(n598), .A1(n597), .B0(n596), .Y(n599) );
  AND2X4TS U1093 ( .A(n573), .B(n2420), .Y(n703) );
  XNOR2X4TS U1094 ( .A(n1505), .B(n551), .Y(addWeight_12__add_s[6]) );
  BUFX8TS U1095 ( .A(n2379), .Y(sumOut[211]) );
  CLKBUFX2TS U1096 ( .A(n2014), .Y(n553) );
  AND2X4TS U1097 ( .A(n898), .B(n2403), .Y(n1875) );
  AND2X4TS U1098 ( .A(n1019), .B(n2440), .Y(n1979) );
  AND2X4TS U1099 ( .A(n994), .B(n2434), .Y(n1839) );
  AND2X4TS U1100 ( .A(n1007), .B(n2437), .Y(n1866) );
  AND2X4TS U1101 ( .A(n873), .B(n2397), .Y(n1857) );
  AND2X4TS U1102 ( .A(n921), .B(n2408), .Y(n1894) );
  AND2X4TS U1103 ( .A(n933), .B(n2411), .Y(n1903) );
  AND2X4TS U1104 ( .A(n970), .B(n2428), .Y(n1930) );
  AND2X4TS U1105 ( .A(n909), .B(n2405), .Y(n1998) );
  AND2X4TS U1106 ( .A(n946), .B(n2422), .Y(n1830) );
  AND2X4TS U1107 ( .A(n982), .B(n2431), .Y(n1848) );
  AND2X4TS U1108 ( .A(n958), .B(n2425), .Y(n1921) );
  AND2X4TS U1109 ( .A(n886), .B(n2400), .Y(n1912) );
  OAI2BB1X4TS U1110 ( .A0N(n1560), .A1N(n1559), .B0(n1558), .Y(n1564) );
  NAND2X4TS U1111 ( .A(n570), .B(n1649), .Y(n575) );
  AND2X4TS U1112 ( .A(n386), .B(n2395), .Y(n1821) );
  AND2X4TS U1113 ( .A(n390), .B(n2390), .Y(n1989) );
  AND2X4TS U1114 ( .A(n826), .B(n2388), .Y(n1970) );
  AND2X4TS U1115 ( .A(n800), .B(n2383), .Y(n1950) );
  AND2X4TS U1116 ( .A(n813), .B(n2386), .Y(n1960) );
  AND2X4TS U1117 ( .A(n787), .B(n2371), .Y(n1940) );
  AND2X4TS U1118 ( .A(n850), .B(n2392), .Y(n1885) );
  NAND2X2TS U1119 ( .A(sumOut[209]), .B(n1442), .Y(n1443) );
  OR2X8TS U1120 ( .A(n2447), .B(n1519), .Y(n1524) );
  OAI2BB1X2TS U1121 ( .A0N(n1285), .A1N(n2014), .B0(n1284), .Y(n1289) );
  OAI2BB1X4TS U1122 ( .A0N(n1497), .A1N(n2010), .B0(n1496), .Y(n1500) );
  OR2X4TS U1123 ( .A(sumOut[153]), .B(n1682), .Y(n1817) );
  OAI21X4TS U1124 ( .A0(n694), .A1(n693), .B0(n692), .Y(n1812) );
  NAND2X2TS U1125 ( .A(n2445), .B(n772), .Y(n657) );
  OR2X8TS U1126 ( .A(n772), .B(n2445), .Y(n1607) );
  NAND2X2TS U1127 ( .A(n2418), .B(n763), .Y(n649) );
  OR2X8TS U1128 ( .A(n763), .B(n2418), .Y(n1603) );
  AOI2BB1X1TS U1129 ( .A0N(sumOut[128]), .A1N(n896), .B0(n628), .Y(
        addWeight_16__add_s[0]) );
  NAND3X2TS U1130 ( .A(n1434), .B(n1478), .C(n1481), .Y(n1439) );
  AND2X4TS U1131 ( .A(n1026), .B(n2369), .Y(n1030) );
  OAI2BB1X2TS U1132 ( .A0N(n1541), .A1N(n1542), .B0(n1540), .Y(n1546) );
  OR2X4TS U1133 ( .A(n2396), .B(n1820), .Y(n858) );
  OAI2BB1X4TS U1134 ( .A0N(n1572), .A1N(n2026), .B0(n1571), .Y(n1576) );
  NAND2X1TS U1135 ( .A(n2042), .B(addWeight_30__add_biasesStored[0]), .Y(n309)
         );
  NAND2X1TS U1136 ( .A(n2031), .B(addWeight_22__add_biasesStored[0]), .Y(n229)
         );
  NAND2X1TS U1137 ( .A(n2046), .B(addWeight_21__add_biasesStored[0]), .Y(n219)
         );
  NAND2X1TS U1138 ( .A(n2039), .B(addWeight_24__add_biasesStored[0]), .Y(n249)
         );
  NAND2BXLTS U1139 ( .AN(addWeight_23__add_biasesStored[0]), .B(n2101), .Y(
        n240) );
  NAND2X1TS U1140 ( .A(n2031), .B(addWeight_20__add_biasesStored[0]), .Y(n209)
         );
  AND2X4TS U1141 ( .A(n1568), .B(n1567), .Y(n1569) );
  OAI2BB1X4TS U1142 ( .A0N(n1274), .A1N(n2014), .B0(n1273), .Y(n1278) );
  OAI2BB1X4TS U1143 ( .A0N(n1280), .A1N(n2022), .B0(n1279), .Y(n1283) );
  INVX2TS U1144 ( .A(n564), .Y(n603) );
  NAND2BX2TS U1145 ( .AN(n600), .B(n599), .Y(n602) );
  OR2X4TS U1146 ( .A(n2374), .B(n677), .Y(n674) );
  INVX2TS U1147 ( .A(n2150), .Y(n835) );
  INVX2TS U1148 ( .A(n2148), .Y(n822) );
  INVX2TS U1149 ( .A(n2138), .Y(n796) );
  INVX2TS U1150 ( .A(n2144), .Y(n809) );
  INVX2TS U1151 ( .A(n2157), .Y(n783) );
  INVX2TS U1152 ( .A(n2155), .Y(n846) );
  INVX2TS U1153 ( .A(n2140), .Y(n859) );
  NAND2X4TS U1154 ( .A(n558), .B(n1660), .Y(n597) );
  INVX2TS U1155 ( .A(n717), .Y(n1027) );
  INVX2TS U1156 ( .A(n571), .Y(n702) );
  INVX2TS U1157 ( .A(weightsIn[53]), .Y(n572) );
  BUFX3TS U1158 ( .A(weightsIn[120]), .Y(n2138) );
  BUFX3TS U1159 ( .A(weightsIn[95]), .Y(n2140) );
  BUFX3TS U1160 ( .A(weightsIn[115]), .Y(n2144) );
  BUFX3TS U1161 ( .A(weightsIn[110]), .Y(n2148) );
  BUFX3TS U1162 ( .A(weightsIn[105]), .Y(n2150) );
  BUFX3TS U1163 ( .A(weightsIn[100]), .Y(n2155) );
  BUFX3TS U1164 ( .A(weightsIn[150]), .Y(n2157) );
  INVX2TS U1165 ( .A(n1452), .Y(n1454) );
  INVX2TS U1166 ( .A(n1245), .Y(n1268) );
  INVX2TS U1167 ( .A(n1433), .Y(n1435) );
  INVX2TS U1168 ( .A(n579), .Y(n582) );
  NOR2X1TS U1169 ( .A(sumOut[229]), .B(n1437), .Y(n1562) );
  INVX2TS U1170 ( .A(n1471), .Y(n1473) );
  INVX2TS U1171 ( .A(n1250), .Y(n1258) );
  INVX2TS U1172 ( .A(sumOut[222]), .Y(n595) );
  INVX2TS U1173 ( .A(n603), .Y(n594) );
  NAND2X1TS U1174 ( .A(sumOut[222]), .B(n603), .Y(n645) );
  AND2X4TS U1175 ( .A(sumOut[4]), .B(n1529), .Y(n2024) );
  AND2X4TS U1176 ( .A(sumOut[252]), .B(n1040), .Y(n2012) );
  AND2X4TS U1177 ( .A(sumOut[100]), .B(n1475), .Y(n2003) );
  AND2X4TS U1178 ( .A(sumOut[212]), .B(n1456), .Y(n2007) );
  OAI21X2TS U1179 ( .A0(sumOut[211]), .A1(n743), .B0(n1441), .Y(n1450) );
  BUFX4TS U1180 ( .A(weightsIn[60]), .Y(n1461) );
  NOR2X4TS U1181 ( .A(sumOut[221]), .B(n605), .Y(n593) );
  NAND2X4TS U1182 ( .A(sumOut[224]), .B(n2164), .Y(n1596) );
  NAND2X2TS U1183 ( .A(n701), .B(n1648), .Y(n2212) );
  AND2X4TS U1184 ( .A(sumOut[156]), .B(n1110), .Y(n1726) );
  INVX2TS U1185 ( .A(n1036), .Y(n1038) );
  OAI21X2TS U1186 ( .A0(n2443), .A1(n589), .B0(n687), .Y(n694) );
  NOR2X2TS U1187 ( .A(n2023), .B(n1580), .Y(n1572) );
  NOR2X1TS U1188 ( .A(n1556), .B(n1562), .Y(n1479) );
  INVX2TS U1189 ( .A(n1526), .Y(n1527) );
  INVX2TS U1190 ( .A(n1417), .Y(n1419) );
  INVX2TS U1191 ( .A(n1425), .Y(n1427) );
  INVX2TS U1192 ( .A(n791), .Y(n1048) );
  INVX2TS U1193 ( .A(n804), .Y(n1058) );
  INVX2TS U1194 ( .A(n817), .Y(n1068) );
  INVX2TS U1195 ( .A(n830), .Y(n1078) );
  INVX2TS U1196 ( .A(n841), .Y(n1088) );
  INVX2TS U1197 ( .A(n854), .Y(n1098) );
  INVX2TS U1198 ( .A(n865), .Y(n1108) );
  INVX2TS U1199 ( .A(n877), .Y(n1118) );
  INVX2TS U1200 ( .A(n890), .Y(n1128) );
  INVX2TS U1201 ( .A(n901), .Y(n1138) );
  INVX2TS U1202 ( .A(n913), .Y(n1148) );
  INVX2TS U1203 ( .A(n925), .Y(n1158) );
  INVX2TS U1204 ( .A(n937), .Y(n1168) );
  INVX2TS U1205 ( .A(n950), .Y(n1178) );
  INVX2TS U1206 ( .A(n962), .Y(n1188) );
  INVX2TS U1207 ( .A(n974), .Y(n1198) );
  INVX2TS U1208 ( .A(n986), .Y(n1208) );
  INVX2TS U1209 ( .A(n998), .Y(n1218) );
  INVX2TS U1210 ( .A(n1011), .Y(n1228) );
  INVX2TS U1211 ( .A(n1023), .Y(n1238) );
  INVX2TS U1212 ( .A(weightsIn[138]), .Y(n623) );
  INVX2TS U1213 ( .A(weightsIn[132]), .Y(n742) );
  OR2X4TS U1214 ( .A(sumOut[98]), .B(n750), .Y(n1460) );
  INVX2TS U1215 ( .A(weightsIn[93]), .Y(n872) );
  INVX2TS U1216 ( .A(weightsIn[88]), .Y(n885) );
  INVX2TS U1217 ( .A(weightsIn[78]), .Y(n908) );
  INVX2TS U1218 ( .A(weightsIn[73]), .Y(n920) );
  INVX2TS U1219 ( .A(weightsIn[43]), .Y(n957) );
  INVX2TS U1220 ( .A(weightsIn[33]), .Y(n981) );
  INVX2TS U1221 ( .A(weightsIn[28]), .Y(n993) );
  INVX2TS U1222 ( .A(weightsIn[18]), .Y(n1018) );
  INVX2TS U1223 ( .A(n785), .Y(n1939) );
  INVX2TS U1224 ( .A(n798), .Y(n1949) );
  INVX2TS U1225 ( .A(n811), .Y(n1959) );
  INVX2TS U1226 ( .A(n824), .Y(n1969) );
  INVX2TS U1227 ( .A(n837), .Y(n1988) );
  INVX2TS U1228 ( .A(n848), .Y(n1884) );
  INVX2TS U1229 ( .A(n861), .Y(n1820) );
  INVX2TS U1230 ( .A(weightsIn[153]), .Y(n786) );
  INVX2TS U1231 ( .A(weightsIn[118]), .Y(n812) );
  INVX2TS U1232 ( .A(weightsIn[113]), .Y(n825) );
  INVX2TS U1233 ( .A(weightsIn[3]), .Y(n711) );
  OR2X4TS U1234 ( .A(sumOut[10]), .B(n659), .Y(n656) );
  OR2X4TS U1235 ( .A(sumOut[90]), .B(n651), .Y(n648) );
  OR2X4TS U1236 ( .A(sumOut[226]), .B(n612), .Y(n609) );
  NOR2X2TS U1237 ( .A(n796), .B(n1945), .Y(n2137) );
  NOR2X2TS U1238 ( .A(n859), .B(n1816), .Y(n2139) );
  NOR2X2TS U1239 ( .A(n809), .B(n1955), .Y(n2143) );
  NOR2X2TS U1240 ( .A(n822), .B(n1965), .Y(n2147) );
  NOR2X2TS U1241 ( .A(n835), .B(n1984), .Y(n2149) );
  NOR2X2TS U1242 ( .A(n846), .B(n1880), .Y(n2154) );
  NOR2X2TS U1243 ( .A(n783), .B(n1935), .Y(n2156) );
  NAND3X2TS U1244 ( .A(n1560), .B(n1479), .C(n1480), .Y(n1434) );
  AND2X4TS U1245 ( .A(n2443), .B(n589), .Y(n690) );
  NAND2X2TS U1246 ( .A(n1444), .B(n2160), .Y(n741) );
  BUFX4TS U1247 ( .A(weightsIn[20]), .Y(n1004) );
  BUFX4TS U1248 ( .A(weightsIn[45]), .Y(n943) );
  BUFX4TS U1249 ( .A(weightsIn[85]), .Y(n883) );
  NOR2BX2TS U1250 ( .AN(n2172), .B(n732), .Y(n2171) );
  NAND2X4TS U1251 ( .A(sumOut[80]), .B(n2142), .Y(n1650) );
  INVX2TS U1252 ( .A(n708), .Y(n2152) );
  INVX2TS U1253 ( .A(n620), .Y(n2151) );
  INVX2TS U1254 ( .A(n722), .Y(n2145) );
  INVX2TS U1255 ( .A(n678), .Y(n676) );
  NAND2X2TS U1256 ( .A(n758), .B(n757), .Y(n1644) );
  NAND2X2TS U1257 ( .A(n766), .B(n765), .Y(n1624) );
  NAND2X2TS U1258 ( .A(n775), .B(n774), .Y(n1634) );
  INVX2TS U1259 ( .A(n869), .Y(n1855) );
  NAND2X2TS U1260 ( .A(n1911), .B(n1910), .Y(n2269) );
  INVX2TS U1261 ( .A(n881), .Y(n1910) );
  NAND2X2TS U1262 ( .A(n1874), .B(n1873), .Y(n2229) );
  INVX2TS U1263 ( .A(n894), .Y(n1873) );
  INVX2TS U1264 ( .A(n905), .Y(n1996) );
  INVX2TS U1265 ( .A(n917), .Y(n1892) );
  NAND2X2TS U1266 ( .A(n1902), .B(n1901), .Y(n2214) );
  INVX2TS U1267 ( .A(n929), .Y(n1901) );
  NAND2X2TS U1268 ( .A(n1829), .B(n1828), .Y(n2204) );
  INVX2TS U1269 ( .A(n941), .Y(n1828) );
  NAND2X2TS U1270 ( .A(n1920), .B(n1919), .Y(n2199) );
  INVX2TS U1271 ( .A(n954), .Y(n1919) );
  NAND2X2TS U1272 ( .A(n1929), .B(n1928), .Y(n2194) );
  INVX2TS U1273 ( .A(n966), .Y(n1928) );
  NAND2X2TS U1274 ( .A(n1847), .B(n1846), .Y(n2189) );
  INVX2TS U1275 ( .A(n978), .Y(n1846) );
  INVX2TS U1276 ( .A(n990), .Y(n1837) );
  NAND2X2TS U1277 ( .A(n1865), .B(n1864), .Y(n2179) );
  INVX2TS U1278 ( .A(n1002), .Y(n1864) );
  INVX2TS U1279 ( .A(n1015), .Y(n1977) );
  CLKAND2X2TS U1280 ( .A(n1235), .B(n1233), .Y(n1024) );
  CLKAND2X2TS U1281 ( .A(n1225), .B(n1223), .Y(n1012) );
  CLKAND2X2TS U1282 ( .A(n1215), .B(n1213), .Y(n999) );
  CLKAND2X2TS U1283 ( .A(n1205), .B(n1203), .Y(n987) );
  CLKAND2X2TS U1284 ( .A(n1195), .B(n1193), .Y(n975) );
  CLKAND2X2TS U1285 ( .A(n1185), .B(n1183), .Y(n963) );
  CLKAND2X2TS U1286 ( .A(n1165), .B(n1163), .Y(n938) );
  CLKAND2X2TS U1287 ( .A(n1155), .B(n1153), .Y(n926) );
  CLKAND2X2TS U1288 ( .A(n1145), .B(n1143), .Y(n914) );
  CLKAND2X2TS U1289 ( .A(n1135), .B(n1133), .Y(n902) );
  CLKAND2X2TS U1290 ( .A(n1125), .B(n1123), .Y(n891) );
  CLKAND2X2TS U1291 ( .A(n1115), .B(n1113), .Y(n878) );
  CLKAND2X2TS U1292 ( .A(n1265), .B(n1263), .Y(n1246) );
  AOI21X1TS U1293 ( .A0(sumOut[223]), .A1(n605), .B0(n604), .Y(n606) );
  NAND3X2TS U1294 ( .A(n602), .B(n645), .C(n642), .Y(n607) );
  CLKAND2X2TS U1295 ( .A(n1255), .B(n1253), .Y(n1251) );
  XOR2X1TS U1296 ( .A(n663), .B(n1542), .Y(addWeight_1__add_s[4]) );
  XOR2X1TS U1297 ( .A(n655), .B(n1551), .Y(addWeight_11__add_s[4]) );
  INVX2TS U1298 ( .A(n2168), .Y(n2169) );
  INVX2TS U1299 ( .A(n2165), .Y(n2166) );
  INVX2TS U1300 ( .A(n2162), .Y(n2163) );
  INVX2TS U1301 ( .A(n748), .Y(n641) );
  XOR2X1TS U1302 ( .A(n720), .B(n719), .Y(addWeight_31__add_s[3]) );
  AOI21X1TS U1303 ( .A0(n2257), .A1(n2254), .B0(n2253), .Y(n720) );
  XOR2X1TS U1304 ( .A(n707), .B(n706), .Y(addWeight_10__add_s[3]) );
  AOI21X1TS U1305 ( .A0(n2212), .A1(n2209), .B0(n2208), .Y(n707) );
  CLKAND2X2TS U1306 ( .A(n1276), .B(n1275), .Y(n1277) );
  CLKAND2X2TS U1307 ( .A(n1045), .B(n1043), .Y(n792) );
  CLKAND2X2TS U1308 ( .A(n1065), .B(n1063), .Y(n818) );
  CLKAND2X2TS U1309 ( .A(n1075), .B(n1073), .Y(n831) );
  CLKAND2X2TS U1310 ( .A(n1085), .B(n1083), .Y(n842) );
  CLKAND2X2TS U1311 ( .A(n1095), .B(n1093), .Y(n855) );
  CLKAND2X2TS U1312 ( .A(n1574), .B(n1573), .Y(n1575) );
  CLKAND2X2TS U1313 ( .A(n1493), .B(n1492), .Y(n1494) );
  CLKAND2X2TS U1314 ( .A(n1487), .B(n1486), .Y(n1488) );
  CLKAND2X2TS U1315 ( .A(n1481), .B(n1480), .Y(n1482) );
  INVX2TS U1316 ( .A(n420), .Y(n588) );
  INVX2TS U1317 ( .A(n572), .Y(n573) );
  INVX2TS U1318 ( .A(n623), .Y(n560) );
  NAND2X2TS U1319 ( .A(sumOut[248]), .B(n556), .Y(n608) );
  INVX2TS U1320 ( .A(n612), .Y(n757) );
  INVX2TS U1321 ( .A(n651), .Y(n765) );
  INVX2TS U1322 ( .A(n659), .Y(n774) );
  INVX2TS U1323 ( .A(n750), .Y(n1459) );
  NAND2X1TS U1324 ( .A(n2382), .B(n2146), .Y(n722) );
  NAND2X2TS U1325 ( .A(sumOut[0]), .B(n2153), .Y(n1713) );
  NAND2X1TS U1326 ( .A(sumOut[0]), .B(n2153), .Y(n708) );
  INVX2TS U1327 ( .A(n686), .Y(n589) );
  INVX2TS U1328 ( .A(n2142), .Y(n568) );
  INVX2TS U1329 ( .A(n2385), .Y(n1945) );
  INVX2TS U1330 ( .A(sumOut[152]), .Y(n1816) );
  INVX2TS U1331 ( .A(sumOut[184]), .Y(n1955) );
  INVX2TS U1332 ( .A(sumOut[176]), .Y(n1965) );
  INVX2TS U1333 ( .A(sumOut[168]), .Y(n1984) );
  INVX2TS U1334 ( .A(n2394), .Y(n1880) );
  INVX2TS U1335 ( .A(sumOut[240]), .Y(n1935) );
  INVX2TS U1336 ( .A(sumOut[10]), .Y(n775) );
  INVX2TS U1337 ( .A(sumOut[90]), .Y(n766) );
  INVX2TS U1338 ( .A(sumOut[98]), .Y(n749) );
  INVX2TS U1339 ( .A(sumOut[226]), .Y(n758) );
  INVX2TS U1340 ( .A(sumOut[26]), .Y(n1978) );
  INVX2TS U1341 ( .A(sumOut[34]), .Y(n1865) );
  INVX2TS U1342 ( .A(sumOut[42]), .Y(n1838) );
  INVX2TS U1343 ( .A(sumOut[50]), .Y(n1847) );
  INVX2TS U1344 ( .A(sumOut[58]), .Y(n1929) );
  INVX2TS U1345 ( .A(sumOut[66]), .Y(n1920) );
  INVX2TS U1346 ( .A(sumOut[74]), .Y(n1829) );
  INVX2TS U1347 ( .A(sumOut[106]), .Y(n1902) );
  INVX2TS U1348 ( .A(sumOut[114]), .Y(n1893) );
  INVX2TS U1349 ( .A(sumOut[122]), .Y(n1997) );
  INVX2TS U1350 ( .A(sumOut[130]), .Y(n1874) );
  INVX2TS U1351 ( .A(sumOut[138]), .Y(n1911) );
  INVX2TS U1352 ( .A(sumOut[146]), .Y(n1856) );
  BUFX4TS U1353 ( .A(weightsIn[51]), .Y(n554) );
  BUFX4TS U1354 ( .A(weightsIn[156]), .Y(n555) );
  INVX2TS U1355 ( .A(weightsIn[139]), .Y(n564) );
  NOR2X4TS U1356 ( .A(sumOut[220]), .B(n605), .Y(n617) );
  BUFX4TS U1357 ( .A(n2378), .Y(sumOut[219]) );
  OR2X4TS U1358 ( .A(sumOut[218]), .B(n559), .Y(n557) );
  OAI21X4TS U1359 ( .A0(sumOut[219]), .A1(n560), .B0(n557), .Y(n598) );
  OR2X8TS U1360 ( .A(sumOut[217]), .B(n396), .Y(n1660) );
  NAND2BX4TS U1361 ( .AN(n2378), .B(n623), .Y(n561) );
  AND2X4TS U1362 ( .A(n560), .B(n2378), .Y(n622) );
  AOI21X4TS U1363 ( .A0(n2263), .A1(n561), .B0(n622), .Y(n596) );
  INVX2TS U1364 ( .A(n618), .Y(n562) );
  NOR2BX2TS U1365 ( .AN(n601), .B(n593), .Y(n565) );
  XOR2X4TS U1366 ( .A(n566), .B(n565), .Y(addWeight_27__add_s[5]) );
  BUFX3TS U1367 ( .A(n2420), .Y(sumOut[83]) );
  CLKINVX1TS U1368 ( .A(weightsIn[52]), .Y(n571) );
  OR2X4TS U1369 ( .A(n2421), .B(n702), .Y(n567) );
  OAI21X4TS U1370 ( .A0(sumOut[83]), .A1(n573), .B0(n567), .Y(n576) );
  NAND2X4TS U1371 ( .A(sumOut[81]), .B(n554), .Y(n569) );
  NAND2X4TS U1372 ( .A(n1650), .B(n569), .Y(n570) );
  OR2X8TS U1373 ( .A(sumOut[81]), .B(n554), .Y(n1649) );
  AOI21X4TS U1374 ( .A0(n704), .A1(n2208), .B0(n703), .Y(n574) );
  OAI21X4TS U1375 ( .A0(n576), .A1(n575), .B0(n574), .Y(n2022) );
  INVX2TS U1376 ( .A(weightsIn[54]), .Y(n577) );
  INVX2TS U1377 ( .A(n577), .Y(n584) );
  NOR2X4TS U1378 ( .A(sumOut[84]), .B(n584), .Y(n2019) );
  NOR2X2TS U1379 ( .A(sumOut[85]), .B(n584), .Y(n1293) );
  AND2X4TS U1380 ( .A(sumOut[85]), .B(n579), .Y(n1292) );
  NOR2X4TS U1381 ( .A(n1292), .B(n2020), .Y(n1279) );
  AOI21X2TS U1382 ( .A0(n2022), .A1(n581), .B0(n580), .Y(n586) );
  NOR2BX1TS U1383 ( .AN(n582), .B(sumOut[87]), .Y(n583) );
  AOI21X1TS U1384 ( .A0(sumOut[87]), .A1(n584), .B0(n583), .Y(n585) );
  XNOR2X1TS U1385 ( .A(n586), .B(n585), .Y(addWeight_10__add_s[7]) );
  NAND2X4TS U1386 ( .A(sumOut[16]), .B(n2159), .Y(n688) );
  BUFX6TS U1387 ( .A(n688), .Y(n1612) );
  INVX4TS U1388 ( .A(n1612), .Y(n2158) );
  NAND2X1TS U1389 ( .A(sumOut[17]), .B(n364), .Y(n1610) );
  OR2X2TS U1390 ( .A(sumOut[18]), .B(n588), .Y(n2294) );
  AND2X8TS U1391 ( .A(sumOut[18]), .B(n588), .Y(n2293) );
  AOI21X4TS U1392 ( .A0(n2297), .A1(n2294), .B0(n462), .Y(n592) );
  INVX2TS U1393 ( .A(n690), .Y(n590) );
  NAND2BX4TS U1394 ( .AN(n2443), .B(n686), .Y(n691) );
  NAND2X1TS U1395 ( .A(n590), .B(n691), .Y(n591) );
  XOR2X4TS U1396 ( .A(n592), .B(n591), .Y(addWeight_2__add_s[3]) );
  XOR2X4TS U1397 ( .A(n607), .B(n606), .Y(addWeight_27__add_s[7]) );
  BUFX3TS U1398 ( .A(n2377), .Y(sumOut[227]) );
  OAI21X4TS U1399 ( .A0(sumOut[227]), .A1(n392), .B0(n609), .Y(n615) );
  NAND2X4TS U1400 ( .A(n610), .B(n1596), .Y(n611) );
  AND2X8TS U1401 ( .A(sumOut[226]), .B(n612), .Y(n1643) );
  AND2X4TS U1402 ( .A(n394), .B(n2377), .Y(n759) );
  AOI21X4TS U1403 ( .A0(n1643), .A1(n760), .B0(n759), .Y(n613) );
  OAI21X4TS U1404 ( .A0(n615), .A1(n614), .B0(n613), .Y(n1560) );
  INVX2TS U1405 ( .A(weightsIn[144]), .Y(n1432) );
  XOR2XLTS U1406 ( .A(n1560), .B(n616), .Y(addWeight_28__add_s[4]) );
  BUFX3TS U1407 ( .A(n2446), .Y(sumOut[8]) );
  BUFX3TS U1408 ( .A(n2395), .Y(sumOut[155]) );
  BUFX3TS U1409 ( .A(n2390), .Y(sumOut[171]) );
  BUFX3TS U1410 ( .A(n2388), .Y(sumOut[179]) );
  BUFX3TS U1411 ( .A(n2383), .Y(sumOut[195]) );
  BUFX3TS U1412 ( .A(n2386), .Y(sumOut[187]) );
  BUFX3TS U1413 ( .A(n2371), .Y(sumOut[243]) );
  BUFX3TS U1414 ( .A(n2392), .Y(sumOut[163]) );
  BUFX3TS U1415 ( .A(n2369), .Y(sumOut[251]) );
  NOR2X1TS U1416 ( .A(n618), .B(n617), .Y(n619) );
  XOR2XLTS U1417 ( .A(n599), .B(n619), .Y(addWeight_27__add_s[4]) );
  NAND2X2TS U1418 ( .A(sumOut[216]), .B(n367), .Y(n620) );
  NAND2X2TS U1419 ( .A(n1660), .B(n2151), .Y(n621) );
  NAND2X1TS U1420 ( .A(sumOut[217]), .B(n396), .Y(n1659) );
  NAND2X2TS U1421 ( .A(n621), .B(n1659), .Y(n2267) );
  OR2X2TS U1422 ( .A(sumOut[218]), .B(n559), .Y(n2264) );
  INVX2TS U1423 ( .A(n622), .Y(n625) );
  XOR2X1TS U1424 ( .A(n627), .B(n626), .Y(addWeight_27__add_s[3]) );
  BUFX3TS U1425 ( .A(n2403), .Y(sumOut[131]) );
  BUFX3TS U1426 ( .A(n2440), .Y(sumOut[27]) );
  BUFX3TS U1427 ( .A(n2434), .Y(sumOut[43]) );
  BUFX3TS U1428 ( .A(n2437), .Y(sumOut[35]) );
  BUFX3TS U1429 ( .A(n2397), .Y(sumOut[147]) );
  BUFX3TS U1430 ( .A(n2408), .Y(sumOut[115]) );
  BUFX3TS U1431 ( .A(n2411), .Y(sumOut[107]) );
  BUFX3TS U1432 ( .A(n2428), .Y(sumOut[59]) );
  BUFX3TS U1433 ( .A(n2405), .Y(sumOut[123]) );
  BUFX3TS U1434 ( .A(n2422), .Y(sumOut[75]) );
  BUFX3TS U1435 ( .A(n2431), .Y(sumOut[51]) );
  BUFX3TS U1436 ( .A(n2425), .Y(sumOut[67]) );
  BUFX3TS U1437 ( .A(n2400), .Y(sumOut[139]) );
  INVX2TS U1438 ( .A(n1872), .Y(n628) );
  NAND2X4TS U1439 ( .A(sumOut[24]), .B(n1017), .Y(n1976) );
  INVX2TS U1440 ( .A(n1976), .Y(n629) );
  NAND2X4TS U1441 ( .A(sumOut[40]), .B(n992), .Y(n1836) );
  INVX2TS U1442 ( .A(n1836), .Y(n630) );
  NAND2X4TS U1443 ( .A(sumOut[32]), .B(n1004), .Y(n1863) );
  INVX2TS U1444 ( .A(n1863), .Y(n631) );
  NAND2X4TS U1445 ( .A(sumOut[144]), .B(n871), .Y(n1854) );
  INVX2TS U1446 ( .A(n1854), .Y(n632) );
  NAND2X4TS U1447 ( .A(sumOut[112]), .B(n919), .Y(n1891) );
  INVX2TS U1448 ( .A(n1891), .Y(n633) );
  NAND2X4TS U1449 ( .A(sumOut[104]), .B(n931), .Y(n1900) );
  INVX2TS U1450 ( .A(n1900), .Y(n634) );
  NAND2X4TS U1451 ( .A(sumOut[56]), .B(n968), .Y(n1927) );
  INVX2TS U1452 ( .A(n1927), .Y(n635) );
  NAND2X4TS U1453 ( .A(sumOut[120]), .B(n907), .Y(n1995) );
  INVX2TS U1454 ( .A(n1995), .Y(n636) );
  NAND2X4TS U1455 ( .A(sumOut[72]), .B(n943), .Y(n1827) );
  INVX2TS U1456 ( .A(n1827), .Y(n637) );
  NAND2X4TS U1457 ( .A(sumOut[48]), .B(n980), .Y(n1845) );
  INVX2TS U1458 ( .A(n1845), .Y(n638) );
  NAND2X4TS U1459 ( .A(sumOut[64]), .B(n956), .Y(n1918) );
  INVX2TS U1460 ( .A(n1918), .Y(n639) );
  NAND2X4TS U1461 ( .A(sumOut[136]), .B(n883), .Y(n1909) );
  INVX2TS U1462 ( .A(n1909), .Y(n640) );
  NAND2X4TS U1463 ( .A(sumOut[96]), .B(n1461), .Y(n748) );
  AOI2BB1X2TS U1464 ( .A0N(sumOut[96]), .A1N(n1461), .B0(n641), .Y(
        addWeight_12__add_s[0]) );
  BUFX3TS U1465 ( .A(n2444), .Y(sumOut[11]) );
  BUFX3TS U1466 ( .A(n2417), .Y(sumOut[91]) );
  AND2X2TS U1467 ( .A(n645), .B(n644), .Y(n646) );
  INVX2TS U1468 ( .A(weightsIn[59]), .Y(n1424) );
  AND2X6TS U1469 ( .A(sumOut[92]), .B(n1429), .Y(n1548) );
  NOR2X4TS U1470 ( .A(sumOut[92]), .B(n1429), .Y(n1547) );
  OAI21X4TS U1471 ( .A0(sumOut[91]), .A1(n380), .B0(n648), .Y(n654) );
  NAND2X2TS U1472 ( .A(n2419), .B(n2167), .Y(n1604) );
  NAND2X2TS U1473 ( .A(n649), .B(n1604), .Y(n650) );
  NAND2X4TS U1474 ( .A(n650), .B(n1603), .Y(n653) );
  AND2X8TS U1475 ( .A(sumOut[90]), .B(n651), .Y(n1623) );
  AND2X4TS U1476 ( .A(n382), .B(n2417), .Y(n767) );
  AOI21X4TS U1477 ( .A0(n1623), .A1(n768), .B0(n767), .Y(n652) );
  OAI21X4TS U1478 ( .A0(n654), .A1(n653), .B0(n652), .Y(n1551) );
  INVX2TS U1479 ( .A(weightsIn[9]), .Y(n1416) );
  AND2X6TS U1480 ( .A(sumOut[12]), .B(n1421), .Y(n1539) );
  OAI21X4TS U1481 ( .A0(sumOut[11]), .A1(n376), .B0(n656), .Y(n662) );
  NAND2X2TS U1482 ( .A(n2446), .B(n2170), .Y(n1608) );
  NAND2X4TS U1483 ( .A(n658), .B(n1607), .Y(n661) );
  AND2X8TS U1484 ( .A(sumOut[10]), .B(n659), .Y(n1633) );
  AND2X4TS U1485 ( .A(n378), .B(n2444), .Y(n776) );
  AOI21X4TS U1486 ( .A0(n1633), .A1(n777), .B0(n776), .Y(n660) );
  OAI21X4TS U1487 ( .A0(n662), .A1(n661), .B0(n660), .Y(n1542) );
  INVX2TS U1488 ( .A(weightsIn[127]), .Y(n668) );
  INVX2TS U1489 ( .A(n668), .Y(n725) );
  NAND2X4TS U1490 ( .A(n667), .B(n721), .Y(n670) );
  INVX2TS U1491 ( .A(n1534), .Y(n1536) );
  NOR2X2TS U1492 ( .A(sumOut[204]), .B(n1536), .Y(n2016) );
  AND2X2TS U1493 ( .A(sumOut[205]), .B(n1536), .Y(n1533) );
  OAI21X4TS U1494 ( .A0(sumOut[235]), .A1(n678), .B0(n674), .Y(n681) );
  NAND2X2TS U1495 ( .A(n2375), .B(n733), .Y(n675) );
  NAND2X2TS U1496 ( .A(n2376), .B(n2172), .Y(n1695) );
  OR2X4TS U1497 ( .A(n733), .B(n2375), .Y(n731) );
  NAND2BX4TS U1498 ( .AN(n2373), .B(n676), .Y(n736) );
  AND2X4TS U1499 ( .A(n2373), .B(n678), .Y(n735) );
  AOI21X4TS U1500 ( .A0(n736), .A1(n1614), .B0(n735), .Y(n679) );
  OAI21X4TS U1501 ( .A0(n681), .A1(n680), .B0(n679), .Y(n1811) );
  INVX2TS U1502 ( .A(weightsIn[149]), .Y(n682) );
  NOR2X1TS U1503 ( .A(sumOut[236]), .B(n1245), .Y(n1809) );
  INVX2TS U1504 ( .A(n682), .Y(n1270) );
  AOI21X2TS U1505 ( .A0(n683), .A1(n1811), .B0(n1808), .Y(n685) );
  AND2X4TS U1506 ( .A(sumOut[237]), .B(n1270), .Y(n1244) );
  NOR2X1TS U1507 ( .A(n1243), .B(n1244), .Y(n684) );
  XNOR2X1TS U1508 ( .A(n685), .B(n684), .Y(addWeight_29__add_s[5]) );
  INVX2TS U1509 ( .A(weightsIn[14]), .Y(n695) );
  NOR2X1TS U1510 ( .A(sumOut[20]), .B(n1250), .Y(n1814) );
  CLKINVX1TS U1511 ( .A(n1814), .Y(n697) );
  NAND2X2TS U1512 ( .A(sumOut[17]), .B(n364), .Y(n689) );
  AOI21X4TS U1513 ( .A0(n691), .A1(n2293), .B0(n690), .Y(n692) );
  INVX2TS U1514 ( .A(n695), .Y(n1260) );
  INVX2TS U1515 ( .A(n1813), .Y(n696) );
  AND2X4TS U1516 ( .A(sumOut[21]), .B(n1260), .Y(n1249) );
  NOR2X1TS U1517 ( .A(n1248), .B(n1249), .Y(n698) );
  NAND2X1TS U1518 ( .A(sumOut[81]), .B(n554), .Y(n1648) );
  OR2X2TS U1519 ( .A(n2421), .B(n702), .Y(n2209) );
  INVX2TS U1520 ( .A(n703), .Y(n705) );
  NAND2X1TS U1521 ( .A(n705), .B(n704), .Y(n706) );
  NAND2X2TS U1522 ( .A(n1521), .B(n2152), .Y(n709) );
  NAND2X1TS U1523 ( .A(sumOut[1]), .B(n362), .Y(n1712) );
  NAND2X2TS U1524 ( .A(n709), .B(n1712), .Y(n1622) );
  OR2X2TS U1525 ( .A(sumOut[2]), .B(n710), .Y(n1619) );
  AOI21X4TS U1526 ( .A0(n1622), .A1(n1619), .B0(n1618), .Y(n714) );
  AND2X4TS U1527 ( .A(n1519), .B(n2447), .Y(n1523) );
  INVX2TS U1528 ( .A(n1523), .Y(n712) );
  XOR2X4TS U1529 ( .A(n714), .B(n713), .Y(addWeight_0__add_s[3]) );
  OR2X8TS U1530 ( .A(n2370), .B(n555), .Y(n1667) );
  CLKINVX1TS U1531 ( .A(weightsIn[157]), .Y(n717) );
  OR2X2TS U1532 ( .A(sumOut[250]), .B(n1027), .Y(n2254) );
  AND2X4TS U1533 ( .A(sumOut[250]), .B(weightsIn[157]), .Y(n2253) );
  INVX2TS U1534 ( .A(n1030), .Y(n718) );
  NAND2X1TS U1535 ( .A(n718), .B(n1031), .Y(n719) );
  INVX2TS U1536 ( .A(n2376), .Y(n732) );
  INVX2TS U1537 ( .A(n732), .Y(sumOut[232]) );
  NAND2X4TS U1538 ( .A(n1670), .B(n2145), .Y(n724) );
  NAND2X4TS U1539 ( .A(n724), .B(n1669), .Y(n2237) );
  AOI21X4TS U1540 ( .A0(n2237), .A1(n2234), .B0(n2233), .Y(n730) );
  INVX2TS U1541 ( .A(n726), .Y(n728) );
  XOR2X4TS U1542 ( .A(n730), .B(n729), .Y(addWeight_25__add_s[3]) );
  NAND2X2TS U1543 ( .A(n731), .B(n2171), .Y(n734) );
  NAND2X1TS U1544 ( .A(sumOut[233]), .B(n733), .Y(n1694) );
  NAND2X2TS U1545 ( .A(n734), .B(n1694), .Y(n1617) );
  OR2X2TS U1546 ( .A(n2374), .B(n677), .Y(n1615) );
  AOI21X4TS U1547 ( .A0(n1617), .A1(n1615), .B0(n1614), .Y(n739) );
  INVX2TS U1548 ( .A(n735), .Y(n737) );
  NAND2X1TS U1549 ( .A(n737), .B(n736), .Y(n738) );
  XOR2X4TS U1550 ( .A(n739), .B(n738), .Y(addWeight_29__add_s[3]) );
  OR2X4TS U1551 ( .A(n1442), .B(sumOut[209]), .Y(n1444) );
  INVX2TS U1552 ( .A(n740), .Y(n2160) );
  NAND2X1TS U1553 ( .A(sumOut[209]), .B(n1442), .Y(n1592) );
  OR2X2TS U1554 ( .A(sumOut[210]), .B(n1440), .Y(n1629) );
  AND2X4TS U1555 ( .A(n743), .B(n2379), .Y(n1446) );
  INVX2TS U1556 ( .A(n1446), .Y(n744) );
  AND2X8TS U1557 ( .A(sumOut[98]), .B(n750), .Y(n1638) );
  AOI21X1TS U1558 ( .A0(n1642), .A1(n1639), .B0(n1638), .Y(n754) );
  AND2X4TS U1559 ( .A(n751), .B(n2414), .Y(n1465) );
  INVX2TS U1560 ( .A(n1465), .Y(n752) );
  NAND2X1TS U1561 ( .A(n1466), .B(n752), .Y(n753) );
  NAND2X2TS U1562 ( .A(sumOut[224]), .B(n2164), .Y(n2162) );
  NAND2X1TS U1563 ( .A(sumOut[225]), .B(n755), .Y(n1595) );
  OAI21X4TS U1564 ( .A0(n2162), .A1(n467), .B0(n1595), .Y(n1647) );
  INVX2TS U1565 ( .A(n759), .Y(n761) );
  NAND2X1TS U1566 ( .A(n761), .B(n760), .Y(n762) );
  NAND2X2TS U1567 ( .A(sumOut[88]), .B(n2167), .Y(n2165) );
  OAI21X4TS U1568 ( .A0(n2165), .A1(n764), .B0(n1602), .Y(n1627) );
  AOI21X4TS U1569 ( .A0(n1627), .A1(n1624), .B0(n1623), .Y(n771) );
  INVX2TS U1570 ( .A(n767), .Y(n769) );
  NAND2X4TS U1571 ( .A(sumOut[8]), .B(n2170), .Y(n2168) );
  OAI21X4TS U1572 ( .A0(n2168), .A1(n773), .B0(n1606), .Y(n1637) );
  AOI21X4TS U1573 ( .A0(n1637), .A1(n1634), .B0(n1633), .Y(n780) );
  INVX2TS U1574 ( .A(n776), .Y(n778) );
  INVX2TS U1575 ( .A(weightsIn[154]), .Y(n781) );
  NOR2X1TS U1576 ( .A(sumOut[244]), .B(n791), .Y(n1788) );
  INVX2TS U1577 ( .A(n781), .Y(n1050) );
  NOR2X1TS U1578 ( .A(n1788), .B(n1413), .Y(n1044) );
  CLKINVX1TS U1579 ( .A(weightsIn[152]), .Y(n785) );
  OR2X4TS U1580 ( .A(sumOut[242]), .B(n1939), .Y(n782) );
  OAI21X4TS U1581 ( .A0(sumOut[243]), .A1(n787), .B0(n782), .Y(n790) );
  NAND2BX4TS U1582 ( .AN(n783), .B(sumOut[240]), .Y(n1710) );
  OAI2BB1X4TS U1583 ( .A0N(n1709), .A1N(n2372), .B0(n1710), .Y(n784) );
  NAND2X4TS U1584 ( .A(n784), .B(n1936), .Y(n789) );
  AND2X4TS U1585 ( .A(sumOut[242]), .B(weightsIn[152]), .Y(n2258) );
  AOI21X4TS U1586 ( .A0(n2258), .A1(n1941), .B0(n1940), .Y(n788) );
  OAI21X4TS U1587 ( .A0(n790), .A1(n789), .B0(n788), .Y(n1790) );
  AND2X4TS U1588 ( .A(sumOut[245]), .B(n1050), .Y(n1412) );
  NAND2BX1TS U1589 ( .AN(n1048), .B(sumOut[246]), .Y(n1045) );
  NAND2BX1TS U1590 ( .AN(sumOut[246]), .B(n1048), .Y(n1043) );
  INVX2TS U1591 ( .A(weightsIn[124]), .Y(n794) );
  NOR2X1TS U1592 ( .A(sumOut[196]), .B(n804), .Y(n1792) );
  INVX2TS U1593 ( .A(n794), .Y(n1060) );
  NOR2X1TS U1594 ( .A(n1792), .B(n1407), .Y(n1054) );
  CLKINVX1TS U1595 ( .A(weightsIn[122]), .Y(n798) );
  OR2X4TS U1596 ( .A(sumOut[194]), .B(n1949), .Y(n795) );
  OAI21X4TS U1597 ( .A0(sumOut[195]), .A1(n800), .B0(n795), .Y(n803) );
  NAND2BX4TS U1598 ( .AN(n796), .B(n2385), .Y(n1655) );
  OAI2BB1X4TS U1599 ( .A0N(n1654), .A1N(n2384), .B0(n1655), .Y(n797) );
  NAND2X4TS U1600 ( .A(n797), .B(n1946), .Y(n802) );
  AND2X4TS U1601 ( .A(sumOut[194]), .B(weightsIn[122]), .Y(n2238) );
  AOI21X4TS U1602 ( .A0(n2238), .A1(n1951), .B0(n1950), .Y(n801) );
  OAI21X4TS U1603 ( .A0(n803), .A1(n802), .B0(n801), .Y(n1794) );
  AND2X4TS U1604 ( .A(sumOut[197]), .B(n1060), .Y(n1406) );
  NAND2BX1TS U1605 ( .AN(n1058), .B(sumOut[198]), .Y(n1055) );
  NAND2BX1TS U1606 ( .AN(sumOut[198]), .B(n1058), .Y(n1053) );
  INVX2TS U1607 ( .A(weightsIn[119]), .Y(n807) );
  NOR2X1TS U1608 ( .A(sumOut[188]), .B(n817), .Y(n1801) );
  INVX2TS U1609 ( .A(n807), .Y(n1070) );
  NOR2X1TS U1610 ( .A(n1801), .B(n1401), .Y(n1064) );
  CLKINVX1TS U1611 ( .A(weightsIn[117]), .Y(n811) );
  OR2X4TS U1612 ( .A(sumOut[186]), .B(n1959), .Y(n808) );
  OAI21X4TS U1613 ( .A0(sumOut[187]), .A1(n813), .B0(n808), .Y(n816) );
  NAND2BX4TS U1614 ( .AN(n809), .B(sumOut[184]), .Y(n1705) );
  OAI2BB1X4TS U1615 ( .A0N(n1704), .A1N(n2387), .B0(n1705), .Y(n810) );
  NAND2X4TS U1616 ( .A(n810), .B(n1956), .Y(n815) );
  AND2X4TS U1617 ( .A(sumOut[186]), .B(weightsIn[117]), .Y(n2273) );
  AOI21X4TS U1618 ( .A0(n2273), .A1(n1961), .B0(n1960), .Y(n814) );
  OAI21X4TS U1619 ( .A0(n816), .A1(n815), .B0(n814), .Y(n1803) );
  AND2X4TS U1620 ( .A(sumOut[189]), .B(n1070), .Y(n1400) );
  NAND2BX1TS U1621 ( .AN(n1068), .B(sumOut[190]), .Y(n1065) );
  NAND2BX1TS U1622 ( .AN(sumOut[190]), .B(n1068), .Y(n1063) );
  INVX2TS U1623 ( .A(weightsIn[114]), .Y(n820) );
  NOR2X1TS U1624 ( .A(sumOut[180]), .B(n830), .Y(n1805) );
  INVX2TS U1625 ( .A(n820), .Y(n1080) );
  NOR2X1TS U1626 ( .A(n1805), .B(n1395), .Y(n1074) );
  CLKINVX1TS U1627 ( .A(weightsIn[112]), .Y(n824) );
  OR2X4TS U1628 ( .A(sumOut[178]), .B(n1969), .Y(n821) );
  OAI21X4TS U1629 ( .A0(sumOut[179]), .A1(n826), .B0(n821), .Y(n829) );
  NAND2BX4TS U1630 ( .AN(n822), .B(sumOut[176]), .Y(n1692) );
  OAI2BB1X4TS U1631 ( .A0N(n1691), .A1N(n2389), .B0(n1692), .Y(n823) );
  NAND2X4TS U1632 ( .A(n823), .B(n1966), .Y(n828) );
  AND2X4TS U1633 ( .A(sumOut[178]), .B(weightsIn[112]), .Y(n2288) );
  AOI21X4TS U1634 ( .A0(n2288), .A1(n1971), .B0(n1970), .Y(n827) );
  OAI21X4TS U1635 ( .A0(n829), .A1(n828), .B0(n827), .Y(n1807) );
  AND2X4TS U1636 ( .A(sumOut[181]), .B(n1080), .Y(n1394) );
  NAND2BX1TS U1637 ( .AN(n1078), .B(sumOut[182]), .Y(n1075) );
  NAND2BX1TS U1638 ( .AN(sumOut[182]), .B(n1078), .Y(n1073) );
  INVX2TS U1639 ( .A(weightsIn[109]), .Y(n833) );
  NOR2X1TS U1640 ( .A(sumOut[172]), .B(n841), .Y(n1745) );
  INVX2TS U1641 ( .A(n833), .Y(n1090) );
  NOR2X1TS U1642 ( .A(n1745), .B(n1389), .Y(n1084) );
  CLKINVX1TS U1643 ( .A(weightsIn[107]), .Y(n837) );
  OR2X4TS U1644 ( .A(sumOut[170]), .B(n1988), .Y(n834) );
  OAI21X4TS U1645 ( .A0(sumOut[171]), .A1(n388), .B0(n834), .Y(n840) );
  NAND2BX4TS U1646 ( .AN(n835), .B(sumOut[168]), .Y(n1664) );
  OAI2BB1X4TS U1647 ( .A0N(n1663), .A1N(n2391), .B0(n1664), .Y(n836) );
  NAND2X4TS U1648 ( .A(n836), .B(n1985), .Y(n839) );
  AND2X4TS U1649 ( .A(sumOut[170]), .B(weightsIn[107]), .Y(n2278) );
  AOI21X4TS U1650 ( .A0(n2278), .A1(n1990), .B0(n1989), .Y(n838) );
  OAI21X4TS U1651 ( .A0(n840), .A1(n839), .B0(n838), .Y(n1747) );
  AND2X4TS U1652 ( .A(sumOut[173]), .B(n1090), .Y(n1388) );
  NAND2BX1TS U1653 ( .AN(n1088), .B(sumOut[174]), .Y(n1085) );
  NAND2BX1TS U1654 ( .AN(sumOut[174]), .B(n1088), .Y(n1083) );
  INVX2TS U1655 ( .A(weightsIn[104]), .Y(n844) );
  NOR2X1TS U1656 ( .A(sumOut[164]), .B(n854), .Y(n1741) );
  INVX2TS U1657 ( .A(n844), .Y(n1100) );
  NOR2X1TS U1658 ( .A(n1741), .B(n1383), .Y(n1094) );
  CLKINVX1TS U1659 ( .A(weightsIn[102]), .Y(n848) );
  OR2X4TS U1660 ( .A(sumOut[162]), .B(n1884), .Y(n845) );
  OAI21X4TS U1661 ( .A0(sumOut[163]), .A1(n850), .B0(n845), .Y(n853) );
  NAND2BX4TS U1662 ( .AN(n846), .B(n2394), .Y(n1674) );
  OAI2BB1X4TS U1663 ( .A0N(n1673), .A1N(n2393), .B0(n1674), .Y(n847) );
  NAND2X4TS U1664 ( .A(n847), .B(n1881), .Y(n852) );
  AND2X4TS U1665 ( .A(sumOut[162]), .B(weightsIn[102]), .Y(n2243) );
  AOI21X4TS U1666 ( .A0(n2243), .A1(n1886), .B0(n1885), .Y(n851) );
  OAI21X4TS U1667 ( .A0(n853), .A1(n852), .B0(n851), .Y(n1743) );
  AND2X4TS U1668 ( .A(sumOut[165]), .B(n1100), .Y(n1382) );
  NAND2BX1TS U1669 ( .AN(n1098), .B(sumOut[166]), .Y(n1095) );
  NAND2BX1TS U1670 ( .AN(sumOut[166]), .B(n1098), .Y(n1093) );
  INVX2TS U1671 ( .A(weightsIn[99]), .Y(n857) );
  NOR2X1TS U1672 ( .A(sumOut[156]), .B(n865), .Y(n1727) );
  INVX2TS U1673 ( .A(n857), .Y(n1110) );
  NOR2X1TS U1674 ( .A(n1727), .B(n1377), .Y(n1104) );
  CLKINVX1TS U1675 ( .A(weightsIn[97]), .Y(n861) );
  OAI21X4TS U1676 ( .A0(sumOut[155]), .A1(n384), .B0(n858), .Y(n864) );
  NAND2BX4TS U1677 ( .AN(n859), .B(sumOut[152]), .Y(n1683) );
  AOI21X4TS U1678 ( .A0(n2283), .A1(n1822), .B0(n1821), .Y(n862) );
  OAI21X4TS U1679 ( .A0(n863), .A1(n864), .B0(n862), .Y(n1729) );
  AND2X4TS U1680 ( .A(sumOut[157]), .B(n1110), .Y(n1376) );
  NAND2BX1TS U1681 ( .AN(n1108), .B(sumOut[158]), .Y(n1105) );
  NAND2BX1TS U1682 ( .AN(sumOut[158]), .B(n1108), .Y(n1103) );
  INVX2TS U1683 ( .A(weightsIn[94]), .Y(n868) );
  NOR2X1TS U1684 ( .A(sumOut[148]), .B(n877), .Y(n1765) );
  INVX2TS U1685 ( .A(n868), .Y(n1120) );
  NOR2X1TS U1686 ( .A(n1765), .B(n1371), .Y(n1114) );
  OR2X4TS U1687 ( .A(sumOut[146]), .B(n869), .Y(n870) );
  OAI21X4TS U1688 ( .A0(sumOut[147]), .A1(n873), .B0(n870), .Y(n876) );
  AND2X8TS U1689 ( .A(sumOut[146]), .B(n869), .Y(n2248) );
  AOI21X4TS U1690 ( .A0(n2248), .A1(n1858), .B0(n1857), .Y(n874) );
  OAI21X4TS U1691 ( .A0(n876), .A1(n875), .B0(n874), .Y(n1763) );
  AND2X4TS U1692 ( .A(sumOut[149]), .B(n1120), .Y(n1370) );
  NAND2BX1TS U1693 ( .AN(n1118), .B(sumOut[150]), .Y(n1115) );
  NAND2BX1TS U1694 ( .AN(sumOut[150]), .B(n1118), .Y(n1113) );
  INVX2TS U1695 ( .A(weightsIn[89]), .Y(n880) );
  NOR2X1TS U1696 ( .A(sumOut[140]), .B(n890), .Y(n1779) );
  INVX2TS U1697 ( .A(n880), .Y(n1130) );
  NOR2X1TS U1698 ( .A(n1779), .B(n1365), .Y(n1124) );
  OR2X4TS U1699 ( .A(sumOut[138]), .B(n881), .Y(n882) );
  OAI21X4TS U1700 ( .A0(sumOut[139]), .A1(n886), .B0(n882), .Y(n889) );
  AND2X8TS U1701 ( .A(sumOut[138]), .B(n881), .Y(n2268) );
  AOI21X4TS U1702 ( .A0(n2268), .A1(n1913), .B0(n1912), .Y(n887) );
  OAI21X4TS U1703 ( .A0(n889), .A1(n888), .B0(n887), .Y(n1777) );
  AND2X4TS U1704 ( .A(sumOut[141]), .B(n1130), .Y(n1364) );
  NAND2BX1TS U1705 ( .AN(n1128), .B(sumOut[142]), .Y(n1125) );
  NAND2BX1TS U1706 ( .AN(sumOut[142]), .B(n1128), .Y(n1123) );
  INVX2TS U1707 ( .A(weightsIn[84]), .Y(n893) );
  NOR2X1TS U1708 ( .A(sumOut[132]), .B(n901), .Y(n1760) );
  INVX2TS U1709 ( .A(n893), .Y(n1140) );
  NOR2X1TS U1710 ( .A(n1760), .B(n1359), .Y(n1134) );
  OR2X4TS U1711 ( .A(sumOut[130]), .B(n894), .Y(n895) );
  OAI21X4TS U1712 ( .A0(sumOut[131]), .A1(n898), .B0(n895), .Y(n900) );
  AND2X8TS U1713 ( .A(sumOut[130]), .B(n894), .Y(n2228) );
  AOI21X4TS U1714 ( .A0(n2228), .A1(n1876), .B0(n1875), .Y(n899) );
  AND2X4TS U1715 ( .A(sumOut[133]), .B(n1140), .Y(n1358) );
  NAND2BX1TS U1716 ( .AN(n1138), .B(sumOut[134]), .Y(n1135) );
  NAND2BX1TS U1717 ( .AN(sumOut[134]), .B(n1138), .Y(n1133) );
  INVX2TS U1718 ( .A(weightsIn[79]), .Y(n904) );
  NOR2X1TS U1719 ( .A(sumOut[124]), .B(n913), .Y(n1737) );
  INVX2TS U1720 ( .A(n904), .Y(n1150) );
  NOR2X1TS U1721 ( .A(n1737), .B(n1353), .Y(n1144) );
  OR2X4TS U1722 ( .A(sumOut[122]), .B(n905), .Y(n906) );
  OAI21X4TS U1723 ( .A0(sumOut[123]), .A1(n909), .B0(n906), .Y(n912) );
  AND2X8TS U1724 ( .A(sumOut[122]), .B(n905), .Y(n2223) );
  AOI21X4TS U1725 ( .A0(n2223), .A1(n1999), .B0(n1998), .Y(n910) );
  OAI21X4TS U1726 ( .A0(n912), .A1(n911), .B0(n910), .Y(n1735) );
  AND2X4TS U1727 ( .A(sumOut[125]), .B(n1150), .Y(n1352) );
  NAND2BX1TS U1728 ( .AN(n1148), .B(sumOut[126]), .Y(n1145) );
  NAND2BX1TS U1729 ( .AN(sumOut[126]), .B(n1148), .Y(n1143) );
  INVX2TS U1730 ( .A(weightsIn[74]), .Y(n916) );
  NOR2X1TS U1731 ( .A(sumOut[116]), .B(n925), .Y(n1755) );
  INVX2TS U1732 ( .A(n916), .Y(n1160) );
  NOR2X1TS U1733 ( .A(n1755), .B(n1347), .Y(n1154) );
  OR2X4TS U1734 ( .A(sumOut[114]), .B(n917), .Y(n918) );
  OAI21X4TS U1735 ( .A0(sumOut[115]), .A1(n921), .B0(n918), .Y(n924) );
  AND2X8TS U1736 ( .A(sumOut[114]), .B(n917), .Y(n2218) );
  AOI21X4TS U1737 ( .A0(n2218), .A1(n1895), .B0(n1894), .Y(n922) );
  OAI21X4TS U1738 ( .A0(n924), .A1(n923), .B0(n922), .Y(n1753) );
  AND2X4TS U1739 ( .A(sumOut[117]), .B(n1160), .Y(n1346) );
  NAND2BX1TS U1740 ( .AN(n1158), .B(sumOut[118]), .Y(n1155) );
  NAND2BX1TS U1741 ( .AN(sumOut[118]), .B(n1158), .Y(n1153) );
  INVX2TS U1742 ( .A(weightsIn[69]), .Y(n928) );
  NOR2X1TS U1743 ( .A(sumOut[108]), .B(n937), .Y(n1774) );
  INVX2TS U1744 ( .A(n928), .Y(n1170) );
  NOR2X1TS U1745 ( .A(n1774), .B(n1341), .Y(n1164) );
  OR2X4TS U1746 ( .A(sumOut[106]), .B(n929), .Y(n930) );
  OAI21X4TS U1747 ( .A0(sumOut[107]), .A1(n933), .B0(n930), .Y(n936) );
  AND2X8TS U1748 ( .A(sumOut[106]), .B(n929), .Y(n2213) );
  AOI21X4TS U1749 ( .A0(n2213), .A1(n1904), .B0(n1903), .Y(n934) );
  OAI21X4TS U1750 ( .A0(n936), .A1(n935), .B0(n934), .Y(n1772) );
  AND2X4TS U1751 ( .A(sumOut[109]), .B(n1170), .Y(n1340) );
  NAND2BX1TS U1752 ( .AN(n1168), .B(sumOut[110]), .Y(n1165) );
  NAND2BX1TS U1753 ( .AN(sumOut[110]), .B(n1168), .Y(n1163) );
  INVX2TS U1754 ( .A(weightsIn[49]), .Y(n940) );
  NOR2X1TS U1755 ( .A(sumOut[76]), .B(n950), .Y(n1770) );
  INVX2TS U1756 ( .A(n940), .Y(n1180) );
  NOR2X1TS U1757 ( .A(n1770), .B(n1335), .Y(n1174) );
  OR2X4TS U1758 ( .A(sumOut[74]), .B(n941), .Y(n942) );
  OAI21X4TS U1759 ( .A0(sumOut[75]), .A1(n946), .B0(n942), .Y(n949) );
  AND2X8TS U1760 ( .A(sumOut[74]), .B(n941), .Y(n2203) );
  AOI21X4TS U1761 ( .A0(n2203), .A1(n1831), .B0(n1830), .Y(n947) );
  OAI21X4TS U1762 ( .A0(n949), .A1(n948), .B0(n947), .Y(n1768) );
  AND2X4TS U1763 ( .A(sumOut[77]), .B(n1180), .Y(n1334) );
  NAND2BX1TS U1764 ( .AN(n1178), .B(sumOut[78]), .Y(n1175) );
  NAND2BX1TS U1765 ( .AN(sumOut[78]), .B(n1178), .Y(n1173) );
  INVX2TS U1766 ( .A(weightsIn[44]), .Y(n953) );
  NOR2X1TS U1767 ( .A(sumOut[68]), .B(n962), .Y(n1784) );
  INVX2TS U1768 ( .A(n953), .Y(n1190) );
  NOR2X1TS U1769 ( .A(n1784), .B(n1329), .Y(n1184) );
  OR2X4TS U1770 ( .A(sumOut[66]), .B(n954), .Y(n955) );
  OAI21X4TS U1771 ( .A0(sumOut[67]), .A1(n958), .B0(n955), .Y(n961) );
  AND2X8TS U1772 ( .A(sumOut[66]), .B(n954), .Y(n2198) );
  AOI21X4TS U1773 ( .A0(n2198), .A1(n1922), .B0(n1921), .Y(n959) );
  OAI21X4TS U1774 ( .A0(n961), .A1(n960), .B0(n959), .Y(n1782) );
  AND2X4TS U1775 ( .A(sumOut[69]), .B(n1190), .Y(n1328) );
  NAND2BX1TS U1776 ( .AN(n1188), .B(sumOut[70]), .Y(n1185) );
  NAND2BX1TS U1777 ( .AN(sumOut[70]), .B(n1188), .Y(n1183) );
  INVX2TS U1778 ( .A(weightsIn[39]), .Y(n965) );
  NOR2X1TS U1779 ( .A(sumOut[60]), .B(n974), .Y(n1732) );
  INVX2TS U1780 ( .A(n965), .Y(n1200) );
  NOR2X1TS U1781 ( .A(n1732), .B(n1323), .Y(n1194) );
  OR2X4TS U1782 ( .A(sumOut[58]), .B(n966), .Y(n967) );
  OAI21X4TS U1783 ( .A0(sumOut[59]), .A1(n970), .B0(n967), .Y(n973) );
  AND2X8TS U1784 ( .A(sumOut[58]), .B(n966), .Y(n2193) );
  AOI21X4TS U1785 ( .A0(n2193), .A1(n1931), .B0(n1930), .Y(n971) );
  OAI21X4TS U1786 ( .A0(n973), .A1(n972), .B0(n971), .Y(n1730) );
  AND2X4TS U1787 ( .A(sumOut[61]), .B(n1200), .Y(n1322) );
  NAND2BX1TS U1788 ( .AN(n1198), .B(sumOut[62]), .Y(n1195) );
  NAND2BX1TS U1789 ( .AN(sumOut[62]), .B(n1198), .Y(n1193) );
  INVX2TS U1790 ( .A(weightsIn[34]), .Y(n977) );
  NOR2X1TS U1791 ( .A(sumOut[52]), .B(n986), .Y(n1750) );
  INVX2TS U1792 ( .A(n977), .Y(n1210) );
  NOR2X1TS U1793 ( .A(n1750), .B(n1317), .Y(n1204) );
  OR2X4TS U1794 ( .A(sumOut[50]), .B(n978), .Y(n979) );
  OAI21X4TS U1795 ( .A0(sumOut[51]), .A1(n982), .B0(n979), .Y(n985) );
  AND2X8TS U1796 ( .A(sumOut[50]), .B(n978), .Y(n2188) );
  AOI21X4TS U1797 ( .A0(n2188), .A1(n1849), .B0(n1848), .Y(n983) );
  OAI21X4TS U1798 ( .A0(n985), .A1(n984), .B0(n983), .Y(n1748) );
  AND2X4TS U1799 ( .A(sumOut[53]), .B(n1210), .Y(n1316) );
  NAND2BX1TS U1800 ( .AN(n1208), .B(sumOut[54]), .Y(n1205) );
  NAND2BX1TS U1801 ( .AN(sumOut[54]), .B(n1208), .Y(n1203) );
  INVX2TS U1802 ( .A(weightsIn[29]), .Y(n989) );
  NOR2X1TS U1803 ( .A(sumOut[44]), .B(n998), .Y(n1723) );
  INVX2TS U1804 ( .A(n989), .Y(n1220) );
  NOR2X1TS U1805 ( .A(n1723), .B(n1311), .Y(n1214) );
  OR2X4TS U1806 ( .A(sumOut[42]), .B(n990), .Y(n991) );
  OAI21X4TS U1807 ( .A0(sumOut[43]), .A1(n994), .B0(n991), .Y(n997) );
  AND2X8TS U1808 ( .A(sumOut[42]), .B(n990), .Y(n2183) );
  AOI21X4TS U1809 ( .A0(n2183), .A1(n1840), .B0(n1839), .Y(n995) );
  OAI21X4TS U1810 ( .A0(n997), .A1(n996), .B0(n995), .Y(n1721) );
  AND2X4TS U1811 ( .A(sumOut[45]), .B(n1220), .Y(n1310) );
  NAND2BX1TS U1812 ( .AN(n1218), .B(sumOut[46]), .Y(n1215) );
  NAND2BX1TS U1813 ( .AN(sumOut[46]), .B(n1218), .Y(n1213) );
  INVX2TS U1814 ( .A(weightsIn[24]), .Y(n1001) );
  NOR2X1TS U1815 ( .A(sumOut[36]), .B(n1011), .Y(n1719) );
  INVX2TS U1816 ( .A(n1001), .Y(n1230) );
  NOR2X1TS U1817 ( .A(n1719), .B(n1305), .Y(n1224) );
  OR2X4TS U1818 ( .A(sumOut[34]), .B(n1002), .Y(n1003) );
  OAI21X4TS U1819 ( .A0(sumOut[35]), .A1(n1007), .B0(n1003), .Y(n1010) );
  AND2X8TS U1820 ( .A(sumOut[34]), .B(n1002), .Y(n2178) );
  AOI21X4TS U1821 ( .A0(n2178), .A1(n1867), .B0(n1866), .Y(n1008) );
  OAI21X4TS U1822 ( .A0(n1010), .A1(n1009), .B0(n1008), .Y(n1717) );
  AND2X4TS U1823 ( .A(sumOut[37]), .B(n1230), .Y(n1304) );
  NAND2BX1TS U1824 ( .AN(n1228), .B(sumOut[38]), .Y(n1225) );
  NAND2BX1TS U1825 ( .AN(sumOut[38]), .B(n1228), .Y(n1223) );
  INVX2TS U1826 ( .A(weightsIn[19]), .Y(n1014) );
  NOR2X1TS U1827 ( .A(sumOut[28]), .B(n1023), .Y(n1797) );
  INVX2TS U1828 ( .A(n1014), .Y(n1240) );
  NOR2X1TS U1829 ( .A(n1797), .B(n1299), .Y(n1234) );
  OR2X4TS U1830 ( .A(sumOut[26]), .B(n1015), .Y(n1016) );
  OAI21X4TS U1831 ( .A0(sumOut[27]), .A1(n1019), .B0(n1016), .Y(n1022) );
  AND2X8TS U1832 ( .A(sumOut[26]), .B(n1015), .Y(n2173) );
  AOI21X4TS U1833 ( .A0(n2173), .A1(n1980), .B0(n1979), .Y(n1020) );
  OAI21X4TS U1834 ( .A0(n1022), .A1(n1021), .B0(n1020), .Y(n1795) );
  AND2X4TS U1835 ( .A(sumOut[29]), .B(n1240), .Y(n1298) );
  NAND2BX1TS U1836 ( .AN(n1238), .B(sumOut[30]), .Y(n1235) );
  NAND2BX1TS U1837 ( .AN(sumOut[30]), .B(n1238), .Y(n1233) );
  INVX2TS U1838 ( .A(weightsIn[159]), .Y(n1035) );
  NOR2X2TS U1839 ( .A(sumOut[253]), .B(n1040), .Y(n1287) );
  OR2X4TS U1840 ( .A(sumOut[250]), .B(n1027), .Y(n1028) );
  OAI21X4TS U1841 ( .A0(sumOut[251]), .A1(n1026), .B0(n1028), .Y(n1034) );
  AOI21X4TS U1842 ( .A0(n2253), .A1(n1031), .B0(n1030), .Y(n1032) );
  CLKINVX3TS U1843 ( .A(n1035), .Y(n1036) );
  NAND2BX1TS U1844 ( .AN(sumOut[254]), .B(n1038), .Y(n1275) );
  NAND3X2TS U1845 ( .A(n2014), .B(n1274), .C(n1275), .Y(n1037) );
  AND2X4TS U1846 ( .A(sumOut[253]), .B(n1036), .Y(n1286) );
  NAND2BX1TS U1847 ( .AN(n1038), .B(sumOut[254]), .Y(n1276) );
  NAND3X2TS U1848 ( .A(n1037), .B(n1273), .C(n1276), .Y(n1042) );
  NOR2BX1TS U1849 ( .AN(n1038), .B(sumOut[255]), .Y(n1039) );
  AOI21X2TS U1850 ( .A0(sumOut[255]), .A1(n1040), .B0(n1039), .Y(n1041) );
  XOR2X4TS U1851 ( .A(n1042), .B(n1041), .Y(addWeight_31__add_s[7]) );
  NAND3X2TS U1852 ( .A(n1790), .B(n1044), .C(n1043), .Y(n1047) );
  NAND3X2TS U1853 ( .A(n1047), .B(n1046), .C(n1045), .Y(n1052) );
  NOR2BX1TS U1854 ( .AN(n1048), .B(sumOut[247]), .Y(n1049) );
  AOI21X2TS U1855 ( .A0(sumOut[247]), .A1(n1050), .B0(n1049), .Y(n1051) );
  XOR2X4TS U1856 ( .A(n1052), .B(n1051), .Y(addWeight_30__add_s[7]) );
  NAND3X2TS U1857 ( .A(n1794), .B(n1054), .C(n1053), .Y(n1057) );
  NOR2BX1TS U1858 ( .AN(n1058), .B(sumOut[199]), .Y(n1059) );
  AOI21X2TS U1859 ( .A0(sumOut[199]), .A1(n1060), .B0(n1059), .Y(n1061) );
  XOR2X4TS U1860 ( .A(n1062), .B(n1061), .Y(addWeight_24__add_s[7]) );
  NAND3X2TS U1861 ( .A(n1803), .B(n1064), .C(n1063), .Y(n1067) );
  NAND3X2TS U1862 ( .A(n1067), .B(n1066), .C(n1065), .Y(n1072) );
  NOR2BX1TS U1863 ( .AN(n1068), .B(sumOut[191]), .Y(n1069) );
  AOI21X2TS U1864 ( .A0(sumOut[191]), .A1(n1070), .B0(n1069), .Y(n1071) );
  XOR2X4TS U1865 ( .A(n1072), .B(n1071), .Y(addWeight_23__add_s[7]) );
  NAND3X2TS U1866 ( .A(n1807), .B(n1074), .C(n1073), .Y(n1077) );
  NAND3X2TS U1867 ( .A(n1077), .B(n1076), .C(n1075), .Y(n1082) );
  NOR2BX1TS U1868 ( .AN(n1078), .B(sumOut[183]), .Y(n1079) );
  AOI21X2TS U1869 ( .A0(sumOut[183]), .A1(n1080), .B0(n1079), .Y(n1081) );
  XOR2X4TS U1870 ( .A(n1082), .B(n1081), .Y(addWeight_22__add_s[7]) );
  NAND3X2TS U1871 ( .A(n1747), .B(n1084), .C(n1083), .Y(n1087) );
  NAND3X2TS U1872 ( .A(n1087), .B(n1086), .C(n1085), .Y(n1092) );
  NOR2BX1TS U1873 ( .AN(n1088), .B(sumOut[175]), .Y(n1089) );
  AOI21X2TS U1874 ( .A0(sumOut[175]), .A1(n1090), .B0(n1089), .Y(n1091) );
  XOR2X4TS U1875 ( .A(n1092), .B(n1091), .Y(addWeight_21__add_s[7]) );
  NAND3X2TS U1876 ( .A(n1743), .B(n1094), .C(n1093), .Y(n1097) );
  NOR2BX1TS U1877 ( .AN(n1098), .B(sumOut[167]), .Y(n1099) );
  AOI21X2TS U1878 ( .A0(sumOut[167]), .A1(n1100), .B0(n1099), .Y(n1101) );
  XOR2X4TS U1879 ( .A(n1102), .B(n1101), .Y(addWeight_20__add_s[7]) );
  NAND3X2TS U1880 ( .A(n1729), .B(n1104), .C(n1103), .Y(n1107) );
  NAND3X2TS U1881 ( .A(n1107), .B(n1106), .C(n1105), .Y(n1112) );
  NOR2BX1TS U1882 ( .AN(n1108), .B(sumOut[159]), .Y(n1109) );
  AOI21X2TS U1883 ( .A0(sumOut[159]), .A1(n1110), .B0(n1109), .Y(n1111) );
  XOR2X4TS U1884 ( .A(n1112), .B(n1111), .Y(addWeight_19__add_s[7]) );
  NAND3X2TS U1885 ( .A(n1763), .B(n1114), .C(n1113), .Y(n1117) );
  NAND3X2TS U1886 ( .A(n1117), .B(n1116), .C(n1115), .Y(n1122) );
  NOR2BX1TS U1887 ( .AN(n1118), .B(sumOut[151]), .Y(n1119) );
  AOI21X2TS U1888 ( .A0(sumOut[151]), .A1(n1120), .B0(n1119), .Y(n1121) );
  XOR2X4TS U1889 ( .A(n1122), .B(n1121), .Y(addWeight_18__add_s[7]) );
  NAND3X2TS U1890 ( .A(n1777), .B(n1124), .C(n1123), .Y(n1127) );
  NAND3X2TS U1891 ( .A(n1127), .B(n1126), .C(n1125), .Y(n1132) );
  NOR2BX1TS U1892 ( .AN(n1128), .B(sumOut[143]), .Y(n1129) );
  AOI21X2TS U1893 ( .A0(sumOut[143]), .A1(n1130), .B0(n1129), .Y(n1131) );
  XOR2X4TS U1894 ( .A(n1132), .B(n1131), .Y(addWeight_17__add_s[7]) );
  NAND3X2TS U1895 ( .A(n1758), .B(n1134), .C(n1133), .Y(n1137) );
  NAND3X2TS U1896 ( .A(n1137), .B(n1136), .C(n1135), .Y(n1142) );
  NOR2BX1TS U1897 ( .AN(n1138), .B(sumOut[135]), .Y(n1139) );
  AOI21X2TS U1898 ( .A0(sumOut[135]), .A1(n1140), .B0(n1139), .Y(n1141) );
  XOR2X4TS U1899 ( .A(n1142), .B(n1141), .Y(addWeight_16__add_s[7]) );
  NAND3X2TS U1900 ( .A(n1735), .B(n1144), .C(n1143), .Y(n1147) );
  NAND3X2TS U1901 ( .A(n1147), .B(n1146), .C(n1145), .Y(n1152) );
  NOR2BX1TS U1902 ( .AN(n1148), .B(sumOut[127]), .Y(n1149) );
  AOI21X2TS U1903 ( .A0(sumOut[127]), .A1(n1150), .B0(n1149), .Y(n1151) );
  XOR2X4TS U1904 ( .A(n1152), .B(n1151), .Y(addWeight_15__add_s[7]) );
  NAND3X2TS U1905 ( .A(n1753), .B(n1154), .C(n1153), .Y(n1157) );
  NAND3X2TS U1906 ( .A(n1157), .B(n1156), .C(n1155), .Y(n1162) );
  NOR2BX1TS U1907 ( .AN(n1158), .B(sumOut[119]), .Y(n1159) );
  AOI21X2TS U1908 ( .A0(sumOut[119]), .A1(n1160), .B0(n1159), .Y(n1161) );
  XOR2X4TS U1909 ( .A(n1162), .B(n1161), .Y(addWeight_14__add_s[7]) );
  NAND3X2TS U1910 ( .A(n1772), .B(n1164), .C(n1163), .Y(n1167) );
  NAND3X2TS U1911 ( .A(n1167), .B(n1166), .C(n1165), .Y(n1172) );
  NOR2BX1TS U1912 ( .AN(n1168), .B(sumOut[111]), .Y(n1169) );
  AOI21X2TS U1913 ( .A0(sumOut[111]), .A1(n1170), .B0(n1169), .Y(n1171) );
  XOR2X4TS U1914 ( .A(n1172), .B(n1171), .Y(addWeight_13__add_s[7]) );
  NAND3X2TS U1915 ( .A(n1768), .B(n1174), .C(n1173), .Y(n1177) );
  NAND3X2TS U1916 ( .A(n1177), .B(n1176), .C(n1175), .Y(n1182) );
  NOR2BX1TS U1917 ( .AN(n1178), .B(sumOut[79]), .Y(n1179) );
  AOI21X2TS U1918 ( .A0(sumOut[79]), .A1(n1180), .B0(n1179), .Y(n1181) );
  XOR2X4TS U1919 ( .A(n1182), .B(n1181), .Y(addWeight_9__add_s[7]) );
  NAND3X2TS U1920 ( .A(n1782), .B(n1184), .C(n1183), .Y(n1187) );
  NAND3X2TS U1921 ( .A(n1187), .B(n1186), .C(n1185), .Y(n1192) );
  NOR2BX1TS U1922 ( .AN(n1188), .B(sumOut[71]), .Y(n1189) );
  AOI21X2TS U1923 ( .A0(sumOut[71]), .A1(n1190), .B0(n1189), .Y(n1191) );
  XOR2X4TS U1924 ( .A(n1192), .B(n1191), .Y(addWeight_8__add_s[7]) );
  NAND3X2TS U1925 ( .A(n1730), .B(n1194), .C(n1193), .Y(n1197) );
  NAND3X2TS U1926 ( .A(n1197), .B(n1196), .C(n1195), .Y(n1202) );
  NOR2BX1TS U1927 ( .AN(n1198), .B(sumOut[63]), .Y(n1199) );
  AOI21X2TS U1928 ( .A0(sumOut[63]), .A1(n1200), .B0(n1199), .Y(n1201) );
  XOR2X4TS U1929 ( .A(n1202), .B(n1201), .Y(addWeight_7__add_s[7]) );
  NAND3X2TS U1930 ( .A(n1748), .B(n1204), .C(n1203), .Y(n1207) );
  NAND3X2TS U1931 ( .A(n1207), .B(n1206), .C(n1205), .Y(n1212) );
  NOR2BX1TS U1932 ( .AN(n1208), .B(sumOut[55]), .Y(n1209) );
  AOI21X2TS U1933 ( .A0(sumOut[55]), .A1(n1210), .B0(n1209), .Y(n1211) );
  XOR2X4TS U1934 ( .A(n1212), .B(n1211), .Y(addWeight_6__add_s[7]) );
  NAND3X2TS U1935 ( .A(n1721), .B(n1214), .C(n1213), .Y(n1217) );
  NAND3X2TS U1936 ( .A(n1217), .B(n1216), .C(n1215), .Y(n1222) );
  NOR2BX1TS U1937 ( .AN(n1218), .B(sumOut[47]), .Y(n1219) );
  AOI21X2TS U1938 ( .A0(sumOut[47]), .A1(n1220), .B0(n1219), .Y(n1221) );
  XOR2X4TS U1939 ( .A(n1222), .B(n1221), .Y(addWeight_5__add_s[7]) );
  NAND3X2TS U1940 ( .A(n1717), .B(n1224), .C(n1223), .Y(n1227) );
  NAND3X2TS U1941 ( .A(n1227), .B(n1226), .C(n1225), .Y(n1232) );
  NOR2BX1TS U1942 ( .AN(n1228), .B(sumOut[39]), .Y(n1229) );
  AOI21X2TS U1943 ( .A0(sumOut[39]), .A1(n1230), .B0(n1229), .Y(n1231) );
  XOR2X4TS U1944 ( .A(n1232), .B(n1231), .Y(addWeight_4__add_s[7]) );
  NAND3X2TS U1945 ( .A(n1795), .B(n1234), .C(n1233), .Y(n1237) );
  NAND3X2TS U1946 ( .A(n1237), .B(n1236), .C(n1235), .Y(n1242) );
  NOR2BX1TS U1947 ( .AN(n1238), .B(sumOut[31]), .Y(n1239) );
  AOI21X2TS U1948 ( .A0(sumOut[31]), .A1(n1240), .B0(n1239), .Y(n1241) );
  XOR2X4TS U1949 ( .A(n1242), .B(n1241), .Y(addWeight_3__add_s[7]) );
  NOR2X1TS U1950 ( .A(n1809), .B(n1243), .Y(n1264) );
  NAND2BX1TS U1951 ( .AN(n1268), .B(sumOut[238]), .Y(n1265) );
  NAND2BX1TS U1952 ( .AN(sumOut[238]), .B(n1268), .Y(n1263) );
  NOR2X1TS U1953 ( .A(n1814), .B(n1248), .Y(n1254) );
  NAND2BX1TS U1954 ( .AN(n1258), .B(sumOut[22]), .Y(n1255) );
  NAND2BX1TS U1955 ( .AN(sumOut[22]), .B(n1258), .Y(n1253) );
  NAND3X2TS U1956 ( .A(n1812), .B(n1254), .C(n1253), .Y(n1257) );
  NAND3X2TS U1957 ( .A(n1257), .B(n1256), .C(n1255), .Y(n1262) );
  NOR2BX1TS U1958 ( .AN(n1258), .B(sumOut[23]), .Y(n1259) );
  AOI21X2TS U1959 ( .A0(sumOut[23]), .A1(n1260), .B0(n1259), .Y(n1261) );
  XOR2X4TS U1960 ( .A(n1262), .B(n1261), .Y(addWeight_2__add_s[7]) );
  NAND3X2TS U1961 ( .A(n1811), .B(n1264), .C(n1263), .Y(n1267) );
  NAND3X2TS U1962 ( .A(n1267), .B(n1266), .C(n1265), .Y(n1272) );
  NOR2BX1TS U1963 ( .AN(n1268), .B(sumOut[239]), .Y(n1269) );
  AOI21X2TS U1964 ( .A0(sumOut[239]), .A1(n1270), .B0(n1269), .Y(n1271) );
  XOR2X4TS U1965 ( .A(n1272), .B(n1271), .Y(addWeight_29__add_s[7]) );
  INVX2TS U1966 ( .A(n2012), .Y(n1284) );
  XOR2X4TS U1967 ( .A(n1289), .B(n1288), .Y(addWeight_31__add_s[5]) );
  INVX2TS U1968 ( .A(n2020), .Y(n1290) );
  OAI2BB1X4TS U1969 ( .A0N(n1291), .A1N(n2022), .B0(n1290), .Y(n1295) );
  NOR2X1TS U1970 ( .A(n1293), .B(n1292), .Y(n1294) );
  XOR2X4TS U1971 ( .A(n1295), .B(n1294), .Y(addWeight_10__add_s[5]) );
  CLKINVX1TS U1972 ( .A(n1797), .Y(n1297) );
  INVX2TS U1973 ( .A(n1796), .Y(n1296) );
  NOR2X1TS U1974 ( .A(n1299), .B(n1298), .Y(n1300) );
  XOR2X4TS U1975 ( .A(n1301), .B(n1300), .Y(addWeight_3__add_s[5]) );
  CLKINVX1TS U1976 ( .A(n1719), .Y(n1303) );
  INVX2TS U1977 ( .A(n1718), .Y(n1302) );
  OAI2BB1X4TS U1978 ( .A0N(n1303), .A1N(n1717), .B0(n1302), .Y(n1307) );
  NOR2X1TS U1979 ( .A(n1305), .B(n1304), .Y(n1306) );
  XOR2X4TS U1980 ( .A(n1307), .B(n1306), .Y(addWeight_4__add_s[5]) );
  CLKINVX1TS U1981 ( .A(n1723), .Y(n1309) );
  INVX2TS U1982 ( .A(n1722), .Y(n1308) );
  NOR2X1TS U1983 ( .A(n1311), .B(n1310), .Y(n1312) );
  XOR2X4TS U1984 ( .A(n1313), .B(n1312), .Y(addWeight_5__add_s[5]) );
  CLKINVX1TS U1985 ( .A(n1750), .Y(n1315) );
  INVX2TS U1986 ( .A(n1749), .Y(n1314) );
  NOR2X1TS U1987 ( .A(n1317), .B(n1316), .Y(n1318) );
  XOR2X4TS U1988 ( .A(n1319), .B(n1318), .Y(addWeight_6__add_s[5]) );
  CLKINVX1TS U1989 ( .A(n1732), .Y(n1321) );
  INVX2TS U1990 ( .A(n1731), .Y(n1320) );
  NOR2X1TS U1991 ( .A(n1323), .B(n1322), .Y(n1324) );
  XOR2X4TS U1992 ( .A(n1325), .B(n1324), .Y(addWeight_7__add_s[5]) );
  CLKINVX1TS U1993 ( .A(n1784), .Y(n1327) );
  INVX2TS U1994 ( .A(n1783), .Y(n1326) );
  NOR2X1TS U1995 ( .A(n1329), .B(n1328), .Y(n1330) );
  XOR2X4TS U1996 ( .A(n1331), .B(n1330), .Y(addWeight_8__add_s[5]) );
  CLKINVX1TS U1997 ( .A(n1770), .Y(n1333) );
  INVX2TS U1998 ( .A(n1769), .Y(n1332) );
  NOR2X1TS U1999 ( .A(n1335), .B(n1334), .Y(n1336) );
  XOR2X4TS U2000 ( .A(n1337), .B(n1336), .Y(addWeight_9__add_s[5]) );
  CLKINVX1TS U2001 ( .A(n1774), .Y(n1339) );
  INVX2TS U2002 ( .A(n1773), .Y(n1338) );
  NOR2X1TS U2003 ( .A(n1341), .B(n1340), .Y(n1342) );
  XOR2X4TS U2004 ( .A(n1343), .B(n1342), .Y(addWeight_13__add_s[5]) );
  CLKINVX1TS U2005 ( .A(n1755), .Y(n1345) );
  INVX2TS U2006 ( .A(n1754), .Y(n1344) );
  OAI2BB1X4TS U2007 ( .A0N(n1345), .A1N(n1753), .B0(n1344), .Y(n1349) );
  NOR2X1TS U2008 ( .A(n1347), .B(n1346), .Y(n1348) );
  XOR2X4TS U2009 ( .A(n1349), .B(n1348), .Y(addWeight_14__add_s[5]) );
  CLKINVX1TS U2010 ( .A(n1737), .Y(n1351) );
  INVX2TS U2011 ( .A(n1736), .Y(n1350) );
  NOR2X1TS U2012 ( .A(n1353), .B(n1352), .Y(n1354) );
  XOR2X4TS U2013 ( .A(n1355), .B(n1354), .Y(addWeight_15__add_s[5]) );
  CLKINVX1TS U2014 ( .A(n1760), .Y(n1357) );
  INVX2TS U2015 ( .A(n1759), .Y(n1356) );
  NOR2X1TS U2016 ( .A(n1359), .B(n1358), .Y(n1360) );
  XOR2X4TS U2017 ( .A(n1361), .B(n1360), .Y(addWeight_16__add_s[5]) );
  CLKINVX1TS U2018 ( .A(n1779), .Y(n1363) );
  INVX2TS U2019 ( .A(n1778), .Y(n1362) );
  NOR2X1TS U2020 ( .A(n1365), .B(n1364), .Y(n1366) );
  XOR2X4TS U2021 ( .A(n1367), .B(n1366), .Y(addWeight_17__add_s[5]) );
  CLKINVX1TS U2022 ( .A(n1765), .Y(n1369) );
  INVX2TS U2023 ( .A(n1764), .Y(n1368) );
  NOR2X1TS U2024 ( .A(n1371), .B(n1370), .Y(n1372) );
  XOR2X4TS U2025 ( .A(n1373), .B(n1372), .Y(addWeight_18__add_s[5]) );
  CLKINVX1TS U2026 ( .A(n1727), .Y(n1375) );
  INVX2TS U2027 ( .A(n1726), .Y(n1374) );
  OAI2BB1X4TS U2028 ( .A0N(n1375), .A1N(n1729), .B0(n1374), .Y(n1379) );
  NOR2X1TS U2029 ( .A(n1377), .B(n1376), .Y(n1378) );
  XOR2X4TS U2030 ( .A(n1379), .B(n1378), .Y(addWeight_19__add_s[5]) );
  CLKINVX1TS U2031 ( .A(n1741), .Y(n1381) );
  INVX2TS U2032 ( .A(n1740), .Y(n1380) );
  OAI2BB1X4TS U2033 ( .A0N(n1381), .A1N(n1743), .B0(n1380), .Y(n1385) );
  NOR2X1TS U2034 ( .A(n1383), .B(n1382), .Y(n1384) );
  XOR2X4TS U2035 ( .A(n1385), .B(n1384), .Y(addWeight_20__add_s[5]) );
  CLKINVX1TS U2036 ( .A(n1745), .Y(n1387) );
  INVX2TS U2037 ( .A(n1744), .Y(n1386) );
  NOR2X1TS U2038 ( .A(n1389), .B(n1388), .Y(n1390) );
  XOR2X4TS U2039 ( .A(n1391), .B(n1390), .Y(addWeight_21__add_s[5]) );
  CLKINVX1TS U2040 ( .A(n1805), .Y(n1393) );
  INVX2TS U2041 ( .A(n1804), .Y(n1392) );
  NOR2X1TS U2042 ( .A(n1395), .B(n1394), .Y(n1396) );
  XOR2X4TS U2043 ( .A(n1397), .B(n1396), .Y(addWeight_22__add_s[5]) );
  CLKINVX1TS U2044 ( .A(n1801), .Y(n1399) );
  INVX2TS U2045 ( .A(n1800), .Y(n1398) );
  NOR2X1TS U2046 ( .A(n1401), .B(n1400), .Y(n1402) );
  XOR2X4TS U2047 ( .A(n1403), .B(n1402), .Y(addWeight_23__add_s[5]) );
  CLKINVX1TS U2048 ( .A(n1792), .Y(n1405) );
  INVX2TS U2049 ( .A(n1791), .Y(n1404) );
  NOR2X1TS U2050 ( .A(n1407), .B(n1406), .Y(n1408) );
  XOR2X4TS U2051 ( .A(n1409), .B(n1408), .Y(addWeight_24__add_s[5]) );
  CLKINVX1TS U2052 ( .A(n1788), .Y(n1411) );
  INVX2TS U2053 ( .A(n1787), .Y(n1410) );
  NOR2X1TS U2054 ( .A(n1413), .B(n1412), .Y(n1414) );
  XOR2X4TS U2055 ( .A(n1415), .B(n1414), .Y(addWeight_30__add_s[5]) );
  NOR2X2TS U2056 ( .A(sumOut[13]), .B(n1421), .Y(n1544) );
  NAND2BX1TS U2057 ( .AN(sumOut[14]), .B(n1419), .Y(n1492) );
  NAND3X2TS U2058 ( .A(n1542), .B(n1491), .C(n1492), .Y(n1418) );
  AND2X4TS U2059 ( .A(sumOut[13]), .B(n1417), .Y(n1543) );
  NOR2X2TS U2060 ( .A(n1543), .B(n1539), .Y(n1490) );
  NAND2BX1TS U2061 ( .AN(n1419), .B(sumOut[14]), .Y(n1493) );
  NOR2BX1TS U2062 ( .AN(n1419), .B(sumOut[15]), .Y(n1420) );
  AOI21X2TS U2063 ( .A0(sumOut[15]), .A1(n1421), .B0(n1420), .Y(n1422) );
  XOR2X4TS U2064 ( .A(n1423), .B(n1422), .Y(addWeight_1__add_s[7]) );
  NOR2X2TS U2065 ( .A(sumOut[93]), .B(n1429), .Y(n1553) );
  AND2X4TS U2066 ( .A(sumOut[93]), .B(n1425), .Y(n1552) );
  NOR2X2TS U2067 ( .A(n1552), .B(n1548), .Y(n1484) );
  NAND2BX1TS U2068 ( .AN(n1427), .B(sumOut[94]), .Y(n1487) );
  NOR2BX1TS U2069 ( .AN(n1427), .B(sumOut[95]), .Y(n1428) );
  AOI21X2TS U2070 ( .A0(sumOut[95]), .A1(n1429), .B0(n1428), .Y(n1430) );
  XOR2X4TS U2071 ( .A(n1431), .B(n1430), .Y(addWeight_11__add_s[7]) );
  NAND2BX1TS U2072 ( .AN(n1435), .B(sumOut[230]), .Y(n1481) );
  NOR2BX1TS U2073 ( .AN(n1435), .B(sumOut[231]), .Y(n1436) );
  AOI21X2TS U2074 ( .A0(sumOut[231]), .A1(n1437), .B0(n1436), .Y(n1438) );
  XOR2X4TS U2075 ( .A(n1439), .B(n1438), .Y(addWeight_28__add_s[7]) );
  AOI21X4TS U2076 ( .A0(n1628), .A1(n1447), .B0(n1446), .Y(n1448) );
  OAI21X4TS U2077 ( .A0(n1450), .A1(n1449), .B0(n1448), .Y(n2010) );
  INVX2TS U2078 ( .A(weightsIn[134]), .Y(n1451) );
  NOR2X1TS U2079 ( .A(sumOut[212]), .B(n1452), .Y(n2008) );
  INVX2TS U2080 ( .A(n1451), .Y(n1456) );
  NOR2X1TS U2081 ( .A(n2008), .B(n1515), .Y(n1497) );
  NAND2BX1TS U2082 ( .AN(sumOut[214]), .B(n1454), .Y(n1498) );
  NAND3X2TS U2083 ( .A(n2010), .B(n1497), .C(n1498), .Y(n1453) );
  AND2X4TS U2084 ( .A(sumOut[213]), .B(n1456), .Y(n1514) );
  NOR2BX1TS U2085 ( .AN(n1454), .B(sumOut[215]), .Y(n1455) );
  AOI21X2TS U2086 ( .A0(sumOut[215]), .A1(n1456), .B0(n1455), .Y(n1457) );
  XOR2X4TS U2087 ( .A(n1458), .B(n1457), .Y(addWeight_26__add_s[7]) );
  OAI21X4TS U2088 ( .A0(sumOut[99]), .A1(n751), .B0(n1460), .Y(n1469) );
  NAND2BX4TS U2089 ( .AN(n1462), .B(n2416), .Y(n1600) );
  OAI2BB1X4TS U2090 ( .A0N(n1463), .A1N(n2415), .B0(n1600), .Y(n1464) );
  NAND2X4TS U2091 ( .A(n1464), .B(n1599), .Y(n1468) );
  AOI21X4TS U2092 ( .A0(n1638), .A1(n1466), .B0(n1465), .Y(n1467) );
  OAI21X4TS U2093 ( .A0(n1469), .A1(n1468), .B0(n1467), .Y(n2005) );
  INVX2TS U2094 ( .A(weightsIn[64]), .Y(n1470) );
  NOR2X1TS U2095 ( .A(sumOut[100]), .B(n1471), .Y(n2004) );
  INVX2TS U2096 ( .A(n1470), .Y(n1475) );
  NOR2X2TS U2097 ( .A(sumOut[101]), .B(n1475), .Y(n1509) );
  NOR2X1TS U2098 ( .A(n2004), .B(n1509), .Y(n1502) );
  NAND3X2TS U2099 ( .A(n2005), .B(n1502), .C(n1503), .Y(n1472) );
  AND2X4TS U2100 ( .A(sumOut[101]), .B(n1475), .Y(n1508) );
  NAND3X2TS U2101 ( .A(n1472), .B(n1501), .C(n1504), .Y(n1477) );
  NOR2BX1TS U2102 ( .AN(n1473), .B(sumOut[103]), .Y(n1474) );
  AOI21X2TS U2103 ( .A0(sumOut[103]), .A1(n1475), .B0(n1474), .Y(n1476) );
  XOR2X4TS U2104 ( .A(n1477), .B(n1476), .Y(addWeight_12__add_s[7]) );
  OAI2BB1X2TS U2105 ( .A0N(n1485), .A1N(n1551), .B0(n1484), .Y(n1489) );
  OAI2BB1X2TS U2106 ( .A0N(n1491), .A1N(n1542), .B0(n1490), .Y(n1495) );
  CLKINVX1TS U2107 ( .A(n2004), .Y(n1507) );
  INVX2TS U2108 ( .A(n2003), .Y(n1506) );
  XOR2X4TS U2109 ( .A(n1511), .B(n1510), .Y(addWeight_12__add_s[5]) );
  CLKINVX1TS U2110 ( .A(n2008), .Y(n1513) );
  INVX2TS U2111 ( .A(n2007), .Y(n1512) );
  OAI2BB1X4TS U2112 ( .A0N(n1513), .A1N(n2010), .B0(n1512), .Y(n1517) );
  NOR2X1TS U2113 ( .A(n1515), .B(n1514), .Y(n1516) );
  XOR2X4TS U2114 ( .A(n1517), .B(n1516), .Y(addWeight_26__add_s[5]) );
  INVX2TS U2115 ( .A(weightsIn[4]), .Y(n1525) );
  INVX2TS U2116 ( .A(n1525), .Y(n1529) );
  NOR2X2TS U2117 ( .A(sumOut[5]), .B(n1529), .Y(n1580) );
  OR2X4TS U2118 ( .A(sumOut[2]), .B(n710), .Y(n1518) );
  NAND2X2TS U2119 ( .A(n2448), .B(n362), .Y(n1520) );
  AND2X4TS U2120 ( .A(sumOut[5]), .B(n1526), .Y(n1579) );
  NOR2BX1TS U2121 ( .AN(n1527), .B(sumOut[7]), .Y(n1528) );
  AOI21X2TS U2122 ( .A0(sumOut[7]), .A1(n1529), .B0(n1528), .Y(n1530) );
  XOR2X4TS U2123 ( .A(n1531), .B(n1530), .Y(addWeight_0__add_s[7]) );
  NAND2BX1TS U2124 ( .AN(n359), .B(sumOut[206]), .Y(n1568) );
  NOR2X4TS U2125 ( .A(n1533), .B(n2015), .Y(n1565) );
  NOR2BX1TS U2126 ( .AN(n1534), .B(sumOut[207]), .Y(n1535) );
  INVX2TS U2127 ( .A(n1539), .Y(n1540) );
  XOR2X4TS U2128 ( .A(n1546), .B(n1545), .Y(addWeight_1__add_s[5]) );
  INVX2TS U2129 ( .A(n1548), .Y(n1549) );
  NOR2X1TS U2130 ( .A(n1553), .B(n1552), .Y(n1554) );
  XOR2X4TS U2131 ( .A(n1555), .B(n1554), .Y(addWeight_11__add_s[5]) );
  INVX2TS U2132 ( .A(n1557), .Y(n1558) );
  NOR2X1TS U2133 ( .A(n1562), .B(n1561), .Y(n1563) );
  XOR2X4TS U2134 ( .A(n1564), .B(n1563), .Y(addWeight_28__add_s[5]) );
  XOR2X4TS U2135 ( .A(n1570), .B(n1569), .Y(addWeight_25__add_s[6]) );
  INVX2TS U2136 ( .A(n2024), .Y(n1577) );
  NOR2X1TS U2137 ( .A(n1580), .B(n1579), .Y(n1581) );
  XOR2X4TS U2138 ( .A(n1582), .B(n1581), .Y(addWeight_0__add_s[5]) );
  CLKBUFX2TS U2139 ( .A(clr), .Y(n2081) );
  CLKBUFX2TS U2140 ( .A(n2081), .Y(n1583) );
  CLKBUFX2TS U2141 ( .A(n1583), .Y(n2079) );
  CLKBUFX2TS U2142 ( .A(n2079), .Y(n2027) );
  CLKBUFX2TS U2143 ( .A(n2027), .Y(n2042) );
  NAND2X1TS U2144 ( .A(n2042), .B(addWeight_30__add_biasesStored[7]), .Y(n307)
         );
  CLKBUFX2TS U2145 ( .A(n2027), .Y(n2059) );
  NAND2X1TS U2146 ( .A(n2059), .B(addWeight_29__add_biasesStored[7]), .Y(n297)
         );
  CLKBUFX2TS U2147 ( .A(n1583), .Y(n2028) );
  CLKBUFX2TS U2148 ( .A(n2028), .Y(n2055) );
  NAND2X1TS U2149 ( .A(n2055), .B(addWeight_26__add_biasesStored[7]), .Y(n267)
         );
  CLKBUFX2TS U2150 ( .A(n1583), .Y(n1584) );
  CLKBUFX2TS U2151 ( .A(n1584), .Y(n2033) );
  NAND2X1TS U2152 ( .A(n2033), .B(addWeight_24__add_biasesStored[7]), .Y(n247)
         );
  CLKBUFX2TS U2153 ( .A(n2081), .Y(n2029) );
  CLKBUFX2TS U2154 ( .A(n2029), .Y(n2082) );
  CLKBUFX2TS U2155 ( .A(n2082), .Y(n2032) );
  CLKBUFX2TS U2156 ( .A(n2032), .Y(n2051) );
  NAND2X1TS U2157 ( .A(n2051), .B(addWeight_23__add_biasesStored[7]), .Y(n237)
         );
  CLKBUFX2TS U2158 ( .A(n2082), .Y(n2030) );
  CLKBUFX2TS U2159 ( .A(n2030), .Y(n2047) );
  NAND2X1TS U2160 ( .A(n2047), .B(addWeight_21__add_biasesStored[7]), .Y(n217)
         );
  CLKBUFX2TS U2161 ( .A(n2030), .Y(n2046) );
  NAND2X1TS U2162 ( .A(n2046), .B(addWeight_20__add_biasesStored[7]), .Y(n207)
         );
  CLKBUFX2TS U2163 ( .A(n2030), .Y(n2031) );
  NAND2X1TS U2164 ( .A(n2031), .B(addWeight_19__add_biasesStored[7]), .Y(n197)
         );
  CLKBUFX2TS U2165 ( .A(n2029), .Y(n2045) );
  NAND2X1TS U2166 ( .A(n2045), .B(addWeight_18__add_biasesStored[7]), .Y(n187)
         );
  CLKBUFX2TS U2167 ( .A(n2029), .Y(n2037) );
  NAND2X1TS U2168 ( .A(n2037), .B(addWeight_17__add_biasesStored[7]), .Y(n177)
         );
  CLKBUFX2TS U2169 ( .A(n2032), .Y(n2038) );
  NAND2X1TS U2170 ( .A(n2038), .B(addWeight_16__add_biasesStored[7]), .Y(n167)
         );
  CLKBUFX2TS U2171 ( .A(n2032), .Y(n2039) );
  NAND2X1TS U2172 ( .A(n2039), .B(addWeight_15__add_biasesStored[7]), .Y(n157)
         );
  CLKBUFX2TS U2173 ( .A(n1584), .Y(n2053) );
  NAND2X1TS U2174 ( .A(n2053), .B(addWeight_14__add_biasesStored[7]), .Y(n147)
         );
  CLKBUFX2TS U2175 ( .A(n1584), .Y(n2054) );
  NAND2X1TS U2176 ( .A(n2054), .B(addWeight_13__add_biasesStored[7]), .Y(n137)
         );
  CLKBUFX2TS U2177 ( .A(n2028), .Y(n2040) );
  NAND2X1TS U2178 ( .A(n2040), .B(addWeight_9__add_biasesStored[7]), .Y(n97)
         );
  CLKBUFX2TS U2179 ( .A(n2028), .Y(n2043) );
  NAND2X1TS U2180 ( .A(n2043), .B(addWeight_8__add_biasesStored[7]), .Y(n87)
         );
  CLKBUFX2TS U2181 ( .A(n1583), .Y(n1585) );
  CLKBUFX2TS U2182 ( .A(n1585), .Y(n2034) );
  CLKBUFX2TS U2183 ( .A(n2034), .Y(n2057) );
  NAND2X1TS U2184 ( .A(n2057), .B(addWeight_7__add_biasesStored[7]), .Y(n77)
         );
  CLKBUFX2TS U2185 ( .A(n1585), .Y(n1586) );
  CLKBUFX2TS U2186 ( .A(n1586), .Y(n2072) );
  NAND2X1TS U2187 ( .A(n2072), .B(addWeight_6__add_biasesStored[7]), .Y(n67)
         );
  CLKBUFX2TS U2188 ( .A(n1586), .Y(n2058) );
  NAND2X1TS U2189 ( .A(n2058), .B(addWeight_5__add_biasesStored[7]), .Y(n57)
         );
  CLKBUFX2TS U2190 ( .A(n2027), .Y(n2065) );
  NAND2X1TS U2191 ( .A(n2065), .B(addWeight_4__add_biasesStored[7]), .Y(n47)
         );
  NAND2X1TS U2192 ( .A(n2065), .B(addWeight_3__add_biasesStored[7]), .Y(n37)
         );
  CLKBUFX2TS U2193 ( .A(n1585), .Y(n2035) );
  CLKBUFX2TS U2194 ( .A(n2035), .Y(n2069) );
  NAND2X1TS U2195 ( .A(n2069), .B(addWeight_2__add_biasesStored[7]), .Y(n27)
         );
  CLKBUFX2TS U2196 ( .A(n1584), .Y(n2044) );
  NAND2X1TS U2197 ( .A(n2044), .B(addWeight_12__add_biasesStored[7]), .Y(n127)
         );
  CLKBUFX2TS U2198 ( .A(n2035), .Y(n2060) );
  NAND2X1TS U2199 ( .A(n2060), .B(addWeight_1__add_biasesStored[7]), .Y(n17)
         );
  CLKBUFX2TS U2200 ( .A(n2034), .Y(n2061) );
  NAND2X1TS U2201 ( .A(n2061), .B(addWeight_31__add_biasesStored[7]), .Y(n317)
         );
  CLKBUFX2TS U2202 ( .A(n1585), .Y(n2064) );
  CLKBUFX2TS U2203 ( .A(n2064), .Y(n2071) );
  NAND2X1TS U2204 ( .A(n2071), .B(addWeight_25__add_biasesStored[7]), .Y(n257)
         );
  CLKBUFX2TS U2205 ( .A(n2064), .Y(n2068) );
  NAND2X1TS U2206 ( .A(n2068), .B(addWeight_11__add_biasesStored[7]), .Y(n117)
         );
  CLKBUFX2TS U2207 ( .A(n1586), .Y(n2074) );
  NAND2X1TS U2208 ( .A(n2074), .B(addWeight_0__add_biasesStored[7]), .Y(n7) );
  NAND2X1TS U2209 ( .A(n2061), .B(addWeight_27__add_biasesStored[7]), .Y(n277)
         );
  CLKBUFX2TS U2210 ( .A(n2064), .Y(n2067) );
  NAND2X1TS U2211 ( .A(n2067), .B(addWeight_10__add_biasesStored[7]), .Y(n107)
         );
  CLKBUFX2TS U2212 ( .A(n1586), .Y(n2041) );
  NAND2X1TS U2213 ( .A(n2041), .B(addWeight_28__add_biasesStored[7]), .Y(n287)
         );
  CLKBUFX2TS U2214 ( .A(biasWriteEnable), .Y(n2136) );
  CLKBUFX2TS U2215 ( .A(n2136), .Y(n1590) );
  CLKBUFX2TS U2216 ( .A(n1590), .Y(n2134) );
  CLKBUFX2TS U2217 ( .A(n2134), .Y(n2077) );
  CLKBUFX2TS U2218 ( .A(n2077), .Y(n1587) );
  CLKBUFX2TS U2219 ( .A(n1587), .Y(n2359) );
  CLKBUFX2TS U2220 ( .A(n1587), .Y(n2361) );
  CLKBUFX2TS U2221 ( .A(n1587), .Y(n2363) );
  CLKBUFX2TS U2222 ( .A(n1590), .Y(n2299) );
  CLKBUFX2TS U2223 ( .A(n2299), .Y(n2300) );
  CLKBUFX2TS U2224 ( .A(n2300), .Y(n2367) );
  CLKBUFX2TS U2225 ( .A(n2300), .Y(n2368) );
  CLKBUFX2TS U2226 ( .A(n1587), .Y(n2362) );
  CLKBUFX2TS U2227 ( .A(n2134), .Y(n1588) );
  CLKBUFX2TS U2228 ( .A(n1588), .Y(n2354) );
  CLKBUFX2TS U2229 ( .A(n1588), .Y(n2353) );
  CLKBUFX2TS U2230 ( .A(n1588), .Y(n2352) );
  CLKBUFX2TS U2231 ( .A(n1588), .Y(n2351) );
  CLKBUFX2TS U2232 ( .A(n1590), .Y(n2350) );
  CLKBUFX2TS U2233 ( .A(n2136), .Y(n1591) );
  CLKBUFX2TS U2234 ( .A(n1591), .Y(n2135) );
  CLKBUFX2TS U2235 ( .A(n2135), .Y(n1589) );
  CLKBUFX2TS U2236 ( .A(n1589), .Y(n2345) );
  CLKBUFX2TS U2237 ( .A(n1589), .Y(n2344) );
  CLKBUFX2TS U2238 ( .A(n1589), .Y(n2343) );
  CLKBUFX2TS U2239 ( .A(n1589), .Y(n2341) );
  CLKBUFX2TS U2240 ( .A(n2135), .Y(n2075) );
  CLKBUFX2TS U2241 ( .A(n2075), .Y(n2339) );
  CLKBUFX2TS U2242 ( .A(n2075), .Y(n2338) );
  CLKBUFX2TS U2243 ( .A(n2075), .Y(n2337) );
  CLKBUFX2TS U2244 ( .A(n1591), .Y(n2336) );
  CLKBUFX2TS U2245 ( .A(n1590), .Y(n2358) );
  CLKBUFX2TS U2246 ( .A(n1591), .Y(n2333) );
  CLKBUFX2TS U2247 ( .A(n1591), .Y(n2332) );
  NAND2X1TS U2248 ( .A(n1444), .B(n1592), .Y(n1594) );
  XOR2X1TS U2249 ( .A(n1594), .B(n740), .Y(addWeight_26__add_s[1]) );
  XOR2X1TS U2250 ( .A(n1597), .B(n1596), .Y(addWeight_28__add_s[1]) );
  NAND2X1TS U2251 ( .A(n1599), .B(n1598), .Y(n1601) );
  XOR2X1TS U2252 ( .A(n1601), .B(n1600), .Y(addWeight_12__add_s[1]) );
  NAND2X1TS U2253 ( .A(n1603), .B(n1602), .Y(n1605) );
  XOR2X1TS U2254 ( .A(n1605), .B(n2165), .Y(addWeight_11__add_s[1]) );
  NAND2X1TS U2255 ( .A(n1607), .B(n1606), .Y(n1609) );
  XOR2X1TS U2256 ( .A(n1609), .B(n2168), .Y(addWeight_1__add_s[1]) );
  NAND2X1TS U2257 ( .A(n1611), .B(n1610), .Y(n1613) );
  XOR2X1TS U2258 ( .A(n1613), .B(n1612), .Y(addWeight_2__add_s[1]) );
  NAND2X1TS U2259 ( .A(n332), .B(n1615), .Y(n1616) );
  XNOR2X1TS U2260 ( .A(n1617), .B(n1616), .Y(addWeight_29__add_s[2]) );
  INVX2TS U2261 ( .A(n1618), .Y(n1620) );
  NAND2X1TS U2262 ( .A(n1620), .B(n1619), .Y(n1621) );
  XNOR2X1TS U2263 ( .A(n1622), .B(n1621), .Y(addWeight_0__add_s[2]) );
  INVX2TS U2264 ( .A(n1623), .Y(n1625) );
  NAND2X1TS U2265 ( .A(n1625), .B(n1624), .Y(n1626) );
  XNOR2X1TS U2266 ( .A(n1627), .B(n1626), .Y(addWeight_11__add_s[2]) );
  INVX2TS U2267 ( .A(n1628), .Y(n1630) );
  NAND2X1TS U2268 ( .A(n1630), .B(n1629), .Y(n1631) );
  XNOR2X1TS U2269 ( .A(n1632), .B(n1631), .Y(addWeight_26__add_s[2]) );
  INVX2TS U2270 ( .A(n1633), .Y(n1635) );
  NAND2X1TS U2271 ( .A(n1635), .B(n1634), .Y(n1636) );
  XNOR2X1TS U2272 ( .A(n1637), .B(n1636), .Y(addWeight_1__add_s[2]) );
  INVX2TS U2273 ( .A(n1638), .Y(n1640) );
  NAND2X1TS U2274 ( .A(n1640), .B(n1639), .Y(n1641) );
  XNOR2X1TS U2275 ( .A(n1642), .B(n1641), .Y(addWeight_12__add_s[2]) );
  INVX2TS U2276 ( .A(n1643), .Y(n1645) );
  NAND2X1TS U2277 ( .A(n1645), .B(n1644), .Y(n1646) );
  XNOR2X1TS U2278 ( .A(n1647), .B(n1646), .Y(addWeight_28__add_s[2]) );
  NAND2X1TS U2279 ( .A(n1649), .B(n1648), .Y(n1651) );
  XOR2X1TS U2280 ( .A(n1651), .B(n1650), .Y(addWeight_10__add_s[1]) );
  NAND2X2TS U2281 ( .A(sumOut[105]), .B(n412), .Y(n1899) );
  XOR2X1TS U2282 ( .A(n1653), .B(n1652), .Y(addWeight_13__add_s[1]) );
  NAND2X1TS U2283 ( .A(n1946), .B(n1947), .Y(n1656) );
  XOR2X1TS U2284 ( .A(n1656), .B(n1655), .Y(addWeight_24__add_s[1]) );
  NAND2X2TS U2285 ( .A(sumOut[145]), .B(n419), .Y(n1853) );
  XOR2X1TS U2286 ( .A(n1658), .B(n1657), .Y(addWeight_18__add_s[1]) );
  NAND2X1TS U2287 ( .A(n1660), .B(n1659), .Y(n1662) );
  XOR2X1TS U2288 ( .A(n1662), .B(n1661), .Y(addWeight_27__add_s[1]) );
  NAND2X1TS U2289 ( .A(n1985), .B(n1986), .Y(n1665) );
  XOR2X1TS U2290 ( .A(n1665), .B(n1664), .Y(addWeight_21__add_s[1]) );
  NAND2X1TS U2291 ( .A(n1667), .B(n1666), .Y(n1668) );
  XOR2X1TS U2292 ( .A(n1668), .B(n608), .Y(addWeight_31__add_s[1]) );
  NAND2X1TS U2293 ( .A(n1670), .B(n1669), .Y(n1672) );
  XOR2X1TS U2294 ( .A(n1672), .B(n722), .Y(addWeight_25__add_s[1]) );
  NAND2X1TS U2295 ( .A(n1881), .B(n1882), .Y(n1675) );
  XOR2X1TS U2296 ( .A(n1675), .B(n1674), .Y(addWeight_20__add_s[1]) );
  NAND2X2TS U2297 ( .A(sumOut[73]), .B(n410), .Y(n1826) );
  XOR2X1TS U2298 ( .A(n1677), .B(n1676), .Y(addWeight_9__add_s[1]) );
  NAND2X2TS U2299 ( .A(sumOut[25]), .B(n372), .Y(n1975) );
  XOR2X1TS U2300 ( .A(n1679), .B(n1678), .Y(addWeight_3__add_s[1]) );
  NAND2X2TS U2301 ( .A(sumOut[113]), .B(n414), .Y(n1890) );
  XOR2X1TS U2302 ( .A(n1681), .B(n1680), .Y(addWeight_14__add_s[1]) );
  NAND2X1TS U2303 ( .A(sumOut[153]), .B(n1682), .Y(n1818) );
  NAND2X1TS U2304 ( .A(n1817), .B(n1818), .Y(n1684) );
  XOR2X1TS U2305 ( .A(n1684), .B(n1683), .Y(addWeight_19__add_s[1]) );
  NAND2X2TS U2306 ( .A(sumOut[57]), .B(n406), .Y(n1926) );
  XOR2X1TS U2307 ( .A(n1686), .B(n1685), .Y(addWeight_7__add_s[1]) );
  NAND2X2TS U2308 ( .A(sumOut[33]), .B(n399), .Y(n1862) );
  XOR2X1TS U2309 ( .A(n1688), .B(n1687), .Y(addWeight_4__add_s[1]) );
  NAND2X2TS U2310 ( .A(sumOut[49]), .B(n404), .Y(n1844) );
  XOR2X1TS U2311 ( .A(n1690), .B(n1689), .Y(addWeight_6__add_s[1]) );
  NAND2X1TS U2312 ( .A(n1966), .B(n1967), .Y(n1693) );
  XOR2X1TS U2313 ( .A(n1693), .B(n1692), .Y(addWeight_22__add_s[1]) );
  NAND2X1TS U2314 ( .A(n731), .B(n1694), .Y(n1697) );
  CLKBUFX2TS U2315 ( .A(n1695), .Y(n1696) );
  XOR2X1TS U2316 ( .A(n1697), .B(n1696), .Y(addWeight_29__add_s[1]) );
  NAND2X2TS U2317 ( .A(sumOut[41]), .B(n402), .Y(n1835) );
  XOR2X1TS U2318 ( .A(n1699), .B(n1698), .Y(addWeight_5__add_s[1]) );
  NAND2X2TS U2319 ( .A(sumOut[129]), .B(n369), .Y(n1871) );
  XOR2X1TS U2320 ( .A(n1701), .B(n1700), .Y(addWeight_16__add_s[1]) );
  NAND2X2TS U2321 ( .A(sumOut[137]), .B(n416), .Y(n1908) );
  XOR2X1TS U2322 ( .A(n1703), .B(n1702), .Y(addWeight_17__add_s[1]) );
  NAND2X1TS U2323 ( .A(n1956), .B(n1957), .Y(n1706) );
  XOR2X1TS U2324 ( .A(n1706), .B(n1705), .Y(addWeight_23__add_s[1]) );
  NAND2X2TS U2325 ( .A(sumOut[121]), .B(n374), .Y(n1994) );
  XOR2X1TS U2326 ( .A(n1708), .B(n1707), .Y(addWeight_15__add_s[1]) );
  NAND2X1TS U2327 ( .A(n1936), .B(n1937), .Y(n1711) );
  XOR2X1TS U2328 ( .A(n1711), .B(n1710), .Y(addWeight_30__add_s[1]) );
  NAND2X1TS U2329 ( .A(n1521), .B(n1712), .Y(n1714) );
  XOR2X1TS U2330 ( .A(n1714), .B(n708), .Y(addWeight_0__add_s[1]) );
  NAND2X2TS U2331 ( .A(sumOut[65]), .B(n408), .Y(n1917) );
  XOR2X1TS U2332 ( .A(n1716), .B(n1715), .Y(addWeight_8__add_s[1]) );
  NOR2X1TS U2333 ( .A(n1719), .B(n1718), .Y(n1720) );
  XOR2X1TS U2334 ( .A(n1717), .B(n1720), .Y(addWeight_4__add_s[4]) );
  CLKBUFX2TS U2335 ( .A(n1721), .Y(n1725) );
  NOR2X1TS U2336 ( .A(n1723), .B(n1722), .Y(n1724) );
  XOR2X1TS U2337 ( .A(n1725), .B(n1724), .Y(addWeight_5__add_s[4]) );
  NOR2X1TS U2338 ( .A(n1727), .B(n1726), .Y(n1728) );
  XOR2X1TS U2339 ( .A(n335), .B(n1728), .Y(addWeight_19__add_s[4]) );
  CLKBUFX2TS U2340 ( .A(n1730), .Y(n1734) );
  NOR2X1TS U2341 ( .A(n1732), .B(n1731), .Y(n1733) );
  XOR2X1TS U2342 ( .A(n1734), .B(n1733), .Y(addWeight_7__add_s[4]) );
  CLKBUFX2TS U2343 ( .A(n1735), .Y(n1739) );
  NOR2X1TS U2344 ( .A(n1737), .B(n1736), .Y(n1738) );
  XOR2X1TS U2345 ( .A(n1739), .B(n1738), .Y(addWeight_15__add_s[4]) );
  NOR2X1TS U2346 ( .A(n1741), .B(n1740), .Y(n1742) );
  XOR2X1TS U2347 ( .A(n1743), .B(n1742), .Y(addWeight_20__add_s[4]) );
  NOR2X1TS U2348 ( .A(n1745), .B(n1744), .Y(n1746) );
  XOR2X1TS U2349 ( .A(n1746), .B(n1747), .Y(addWeight_21__add_s[4]) );
  CLKBUFX2TS U2350 ( .A(n1748), .Y(n1752) );
  NOR2X1TS U2351 ( .A(n1750), .B(n1749), .Y(n1751) );
  XOR2X1TS U2352 ( .A(n1752), .B(n1751), .Y(addWeight_6__add_s[4]) );
  CLKBUFX2TS U2353 ( .A(n1753), .Y(n1757) );
  NOR2X1TS U2354 ( .A(n1755), .B(n1754), .Y(n1756) );
  XOR2X1TS U2355 ( .A(n1757), .B(n1756), .Y(addWeight_14__add_s[4]) );
  CLKBUFX2TS U2356 ( .A(n1758), .Y(n1762) );
  NOR2X1TS U2357 ( .A(n1760), .B(n1759), .Y(n1761) );
  XOR2X1TS U2358 ( .A(n1762), .B(n1761), .Y(addWeight_16__add_s[4]) );
  CLKBUFX2TS U2359 ( .A(n1763), .Y(n1767) );
  NOR2X1TS U2360 ( .A(n1765), .B(n1764), .Y(n1766) );
  XOR2X1TS U2361 ( .A(n1767), .B(n1766), .Y(addWeight_18__add_s[4]) );
  NOR2X1TS U2362 ( .A(n1770), .B(n1769), .Y(n1771) );
  XOR2X1TS U2363 ( .A(n1768), .B(n1771), .Y(addWeight_9__add_s[4]) );
  CLKBUFX2TS U2364 ( .A(n1772), .Y(n1776) );
  NOR2X1TS U2365 ( .A(n1774), .B(n1773), .Y(n1775) );
  XOR2X1TS U2366 ( .A(n1776), .B(n1775), .Y(addWeight_13__add_s[4]) );
  CLKBUFX2TS U2367 ( .A(n1777), .Y(n1781) );
  NOR2X1TS U2368 ( .A(n1779), .B(n1778), .Y(n1780) );
  XOR2X1TS U2369 ( .A(n1781), .B(n1780), .Y(addWeight_17__add_s[4]) );
  CLKBUFX2TS U2370 ( .A(n1782), .Y(n1786) );
  NOR2X1TS U2371 ( .A(n1784), .B(n1783), .Y(n1785) );
  XOR2X1TS U2372 ( .A(n1786), .B(n1785), .Y(addWeight_8__add_s[4]) );
  NOR2X1TS U2373 ( .A(n1788), .B(n1787), .Y(n1789) );
  XOR2X1TS U2374 ( .A(n352), .B(n1789), .Y(addWeight_30__add_s[4]) );
  NOR2X1TS U2375 ( .A(n1792), .B(n1791), .Y(n1793) );
  XOR2X1TS U2376 ( .A(n1794), .B(n1793), .Y(addWeight_24__add_s[4]) );
  CLKBUFX2TS U2377 ( .A(n1795), .Y(n1799) );
  NOR2X1TS U2378 ( .A(n1797), .B(n1796), .Y(n1798) );
  XOR2X1TS U2379 ( .A(n1799), .B(n1798), .Y(addWeight_3__add_s[4]) );
  NOR2X1TS U2380 ( .A(n1801), .B(n1800), .Y(n1802) );
  XOR2X1TS U2381 ( .A(n351), .B(n1802), .Y(addWeight_23__add_s[4]) );
  NOR2X1TS U2382 ( .A(n1805), .B(n1804), .Y(n1806) );
  XOR2X1TS U2383 ( .A(n350), .B(n1806), .Y(addWeight_22__add_s[4]) );
  NOR2X1TS U2384 ( .A(n1809), .B(n1808), .Y(n1810) );
  XOR2X1TS U2385 ( .A(n355), .B(n1810), .Y(addWeight_29__add_s[4]) );
  NOR2X1TS U2386 ( .A(n1814), .B(n1813), .Y(n1815) );
  XOR2X1TS U2387 ( .A(n336), .B(n1815), .Y(addWeight_2__add_s[4]) );
  NAND2X2TS U2388 ( .A(n1819), .B(n1818), .Y(n2287) );
  OR2X2TS U2389 ( .A(n2396), .B(n1820), .Y(n2284) );
  AOI21X2TS U2390 ( .A0(n2287), .A1(n2284), .B0(n2283), .Y(n1825) );
  INVX2TS U2391 ( .A(n1821), .Y(n1823) );
  NAND2X1TS U2392 ( .A(n1823), .B(n1822), .Y(n1824) );
  XOR2X1TS U2393 ( .A(n1825), .B(n1824), .Y(addWeight_19__add_s[3]) );
  OAI21X4TS U2394 ( .A0(n1827), .A1(n523), .B0(n1826), .Y(n2207) );
  AOI21X4TS U2395 ( .A0(n2207), .A1(n2204), .B0(n2203), .Y(n1834) );
  INVX2TS U2396 ( .A(n1830), .Y(n1832) );
  NAND2X1TS U2397 ( .A(n1832), .B(n1831), .Y(n1833) );
  XOR2X1TS U2398 ( .A(n1834), .B(n1833), .Y(addWeight_9__add_s[3]) );
  INVX2TS U2399 ( .A(n1839), .Y(n1841) );
  NAND2X1TS U2400 ( .A(n1841), .B(n1840), .Y(n1842) );
  XOR2X1TS U2401 ( .A(n1843), .B(n1842), .Y(addWeight_5__add_s[3]) );
  OAI21X4TS U2402 ( .A0(n1845), .A1(n529), .B0(n1844), .Y(n2192) );
  AOI21X4TS U2403 ( .A0(n2192), .A1(n2189), .B0(n2188), .Y(n1852) );
  INVX2TS U2404 ( .A(n1848), .Y(n1850) );
  NAND2X1TS U2405 ( .A(n1850), .B(n1849), .Y(n1851) );
  XOR2X1TS U2406 ( .A(n1852), .B(n1851), .Y(addWeight_6__add_s[3]) );
  INVX2TS U2407 ( .A(n1857), .Y(n1859) );
  NAND2X1TS U2408 ( .A(n1859), .B(n1858), .Y(n1860) );
  XOR2X1TS U2409 ( .A(n1861), .B(n1860), .Y(addWeight_18__add_s[3]) );
  OAI21X4TS U2410 ( .A0(n1863), .A1(n533), .B0(n1862), .Y(n2182) );
  AOI21X4TS U2411 ( .A0(n2182), .A1(n2179), .B0(n2178), .Y(n1870) );
  INVX2TS U2412 ( .A(n1866), .Y(n1868) );
  NAND2X1TS U2413 ( .A(n1868), .B(n1867), .Y(n1869) );
  XOR2X1TS U2414 ( .A(n1870), .B(n1869), .Y(addWeight_4__add_s[3]) );
  OAI21X4TS U2415 ( .A0(n1872), .A1(n515), .B0(n1871), .Y(n2232) );
  AOI21X4TS U2416 ( .A0(n2232), .A1(n2229), .B0(n2228), .Y(n1879) );
  INVX2TS U2417 ( .A(n1875), .Y(n1877) );
  NAND2X1TS U2418 ( .A(n1877), .B(n1876), .Y(n1878) );
  XOR2X1TS U2419 ( .A(n1879), .B(n1878), .Y(addWeight_16__add_s[3]) );
  NAND2X2TS U2420 ( .A(n1883), .B(n1882), .Y(n2247) );
  OR2X2TS U2421 ( .A(sumOut[162]), .B(n1884), .Y(n2244) );
  INVX2TS U2422 ( .A(n1885), .Y(n1887) );
  NAND2X1TS U2423 ( .A(n1887), .B(n1886), .Y(n1888) );
  XOR2X1TS U2424 ( .A(n1889), .B(n1888), .Y(addWeight_20__add_s[3]) );
  INVX2TS U2425 ( .A(n1894), .Y(n1896) );
  NAND2X1TS U2426 ( .A(n1896), .B(n1895), .Y(n1897) );
  XOR2X1TS U2427 ( .A(n1898), .B(n1897), .Y(addWeight_14__add_s[3]) );
  OAI21X4TS U2428 ( .A0(n1900), .A1(n521), .B0(n1899), .Y(n2217) );
  AOI21X4TS U2429 ( .A0(n2217), .A1(n2214), .B0(n2213), .Y(n1907) );
  INVX2TS U2430 ( .A(n1903), .Y(n1905) );
  NAND2X1TS U2431 ( .A(n1905), .B(n1904), .Y(n1906) );
  XOR2X1TS U2432 ( .A(n1907), .B(n1906), .Y(addWeight_13__add_s[3]) );
  OAI21X4TS U2433 ( .A0(n1909), .A1(n489), .B0(n1908), .Y(n2272) );
  AOI21X4TS U2434 ( .A0(n2272), .A1(n2269), .B0(n2268), .Y(n1916) );
  INVX2TS U2435 ( .A(n1912), .Y(n1914) );
  NAND2X1TS U2436 ( .A(n1914), .B(n1913), .Y(n1915) );
  XOR2X1TS U2437 ( .A(n1916), .B(n1915), .Y(addWeight_17__add_s[3]) );
  OAI21X4TS U2438 ( .A0(n1918), .A1(n525), .B0(n1917), .Y(n2202) );
  AOI21X4TS U2439 ( .A0(n2202), .A1(n2199), .B0(n2198), .Y(n1925) );
  INVX2TS U2440 ( .A(n1921), .Y(n1923) );
  NAND2X1TS U2441 ( .A(n1923), .B(n1922), .Y(n1924) );
  XOR2X1TS U2442 ( .A(n1925), .B(n1924), .Y(addWeight_8__add_s[3]) );
  OAI21X4TS U2443 ( .A0(n1927), .A1(n527), .B0(n1926), .Y(n2197) );
  AOI21X4TS U2444 ( .A0(n2197), .A1(n2194), .B0(n2193), .Y(n1934) );
  INVX2TS U2445 ( .A(n1930), .Y(n1932) );
  NAND2X1TS U2446 ( .A(n1932), .B(n1931), .Y(n1933) );
  XOR2X1TS U2447 ( .A(n1934), .B(n1933), .Y(addWeight_7__add_s[3]) );
  NAND2X2TS U2448 ( .A(n1938), .B(n1937), .Y(n2262) );
  OR2X2TS U2449 ( .A(sumOut[242]), .B(n1939), .Y(n2259) );
  INVX2TS U2450 ( .A(n1940), .Y(n1942) );
  NAND2X1TS U2451 ( .A(n1942), .B(n1941), .Y(n1943) );
  XOR2X1TS U2452 ( .A(n1944), .B(n1943), .Y(addWeight_30__add_s[3]) );
  NAND2X2TS U2453 ( .A(n1948), .B(n1947), .Y(n2242) );
  OR2X2TS U2454 ( .A(sumOut[194]), .B(n1949), .Y(n2239) );
  INVX2TS U2455 ( .A(n1950), .Y(n1952) );
  NAND2X1TS U2456 ( .A(n1952), .B(n1951), .Y(n1953) );
  XOR2X1TS U2457 ( .A(n1954), .B(n1953), .Y(addWeight_24__add_s[3]) );
  NAND2X2TS U2458 ( .A(n1958), .B(n1957), .Y(n2277) );
  OR2X2TS U2459 ( .A(sumOut[186]), .B(n1959), .Y(n2274) );
  INVX2TS U2460 ( .A(n1960), .Y(n1962) );
  NAND2X1TS U2461 ( .A(n1962), .B(n1961), .Y(n1963) );
  XOR2X1TS U2462 ( .A(n1964), .B(n1963), .Y(addWeight_23__add_s[3]) );
  NAND2X2TS U2463 ( .A(n1968), .B(n1967), .Y(n2292) );
  OR2X2TS U2464 ( .A(sumOut[178]), .B(n1969), .Y(n2289) );
  INVX2TS U2465 ( .A(n1970), .Y(n1972) );
  NAND2X1TS U2466 ( .A(n1972), .B(n1971), .Y(n1973) );
  XOR2X1TS U2467 ( .A(n1974), .B(n1973), .Y(addWeight_22__add_s[3]) );
  INVX2TS U2468 ( .A(n1979), .Y(n1981) );
  NAND2X1TS U2469 ( .A(n1981), .B(n1980), .Y(n1982) );
  XOR2X1TS U2470 ( .A(n1983), .B(n1982), .Y(addWeight_3__add_s[3]) );
  NAND2X2TS U2471 ( .A(n1987), .B(n1986), .Y(n2282) );
  OR2X2TS U2472 ( .A(sumOut[170]), .B(n1988), .Y(n2279) );
  INVX2TS U2473 ( .A(n1989), .Y(n1991) );
  NAND2X1TS U2474 ( .A(n1991), .B(n1990), .Y(n1992) );
  XOR2X1TS U2475 ( .A(n1993), .B(n1992), .Y(addWeight_21__add_s[3]) );
  INVX2TS U2476 ( .A(n1998), .Y(n2000) );
  NAND2X1TS U2477 ( .A(n2000), .B(n1999), .Y(n2001) );
  XOR2X1TS U2478 ( .A(n2002), .B(n2001), .Y(addWeight_15__add_s[3]) );
  NOR2X1TS U2479 ( .A(n2004), .B(n2003), .Y(n2006) );
  XOR2X1TS U2480 ( .A(n2006), .B(n2005), .Y(addWeight_12__add_s[4]) );
  NOR2X1TS U2481 ( .A(n2008), .B(n2007), .Y(n2009) );
  XOR2X1TS U2482 ( .A(n2009), .B(n2010), .Y(addWeight_26__add_s[4]) );
  NOR2X1TS U2483 ( .A(n2012), .B(n2011), .Y(n2013) );
  XOR2X1TS U2484 ( .A(n553), .B(n2013), .Y(addWeight_31__add_s[4]) );
  NOR2X1TS U2485 ( .A(n2016), .B(n2015), .Y(n2018) );
  XOR2X1TS U2486 ( .A(n2018), .B(n2017), .Y(addWeight_25__add_s[4]) );
  NOR2X1TS U2487 ( .A(n2020), .B(n2019), .Y(n2021) );
  XOR2X1TS U2488 ( .A(n2021), .B(n2022), .Y(addWeight_10__add_s[4]) );
  NOR2X1TS U2489 ( .A(n2024), .B(n2023), .Y(n2025) );
  XOR2X1TS U2490 ( .A(n2025), .B(n2026), .Y(addWeight_0__add_s[4]) );
  CLKBUFX2TS U2491 ( .A(n2035), .Y(n2070) );
  NAND2X1TS U2492 ( .A(n2070), .B(addWeight_2__add_biasesStored[2]), .Y(n23)
         );
  CLKBUFX2TS U2493 ( .A(n2082), .Y(n2049) );
  NAND2X1TS U2494 ( .A(n2049), .B(addWeight_22__add_biasesStored[7]), .Y(n227)
         );
  NAND2X1TS U2495 ( .A(n2072), .B(addWeight_31__add_biasesStored[1]), .Y(n311)
         );
  NAND2X1TS U2496 ( .A(n2069), .B(addWeight_31__add_biasesStored[0]), .Y(n319)
         );
  CLKBUFX2TS U2497 ( .A(n2027), .Y(n2036) );
  NAND2X1TS U2498 ( .A(n2036), .B(addWeight_30__add_biasesStored[1]), .Y(n301)
         );
  NAND2X1TS U2499 ( .A(n2072), .B(addWeight_29__add_biasesStored[1]), .Y(n291)
         );
  CLKBUFX2TS U2500 ( .A(n2028), .Y(n2056) );
  NAND2X1TS U2501 ( .A(n2056), .B(addWeight_27__add_biasesStored[1]), .Y(n271)
         );
  NAND2X1TS U2502 ( .A(n2040), .B(addWeight_27__add_biasesStored[0]), .Y(n279)
         );
  NAND2X1TS U2503 ( .A(n2054), .B(addWeight_25__add_biasesStored[1]), .Y(n251)
         );
  NAND2X1TS U2504 ( .A(n2033), .B(addWeight_25__add_biasesStored[0]), .Y(n259)
         );
  NAND2X1TS U2505 ( .A(n2039), .B(addWeight_24__add_biasesStored[1]), .Y(n241)
         );
  CLKBUFX2TS U2506 ( .A(n2029), .Y(n2050) );
  NAND2X1TS U2507 ( .A(n2050), .B(addWeight_23__add_biasesStored[1]), .Y(n231)
         );
  NAND2X1TS U2508 ( .A(n2037), .B(addWeight_23__add_biasesStored[0]), .Y(n239)
         );
  CLKBUFX2TS U2509 ( .A(n2030), .Y(n2048) );
  NAND2X1TS U2510 ( .A(n2048), .B(addWeight_22__add_biasesStored[1]), .Y(n221)
         );
  NAND2X1TS U2511 ( .A(n2056), .B(addWeight_21__add_biasesStored[1]), .Y(n211)
         );
  NAND2X1TS U2512 ( .A(n2031), .B(addWeight_20__add_biasesStored[1]), .Y(n201)
         );
  NAND2X1TS U2513 ( .A(n2048), .B(addWeight_19__add_biasesStored[1]), .Y(n191)
         );
  NAND2X1TS U2514 ( .A(n2045), .B(addWeight_19__add_biasesStored[0]), .Y(n199)
         );
  NAND2X1TS U2515 ( .A(n2049), .B(addWeight_18__add_biasesStored[1]), .Y(n181)
         );
  NAND2X1TS U2516 ( .A(n2037), .B(addWeight_18__add_biasesStored[0]), .Y(n189)
         );
  NAND2X1TS U2517 ( .A(n2050), .B(addWeight_17__add_biasesStored[1]), .Y(n171)
         );
  NAND2X1TS U2518 ( .A(n2038), .B(addWeight_17__add_biasesStored[0]), .Y(n179)
         );
  NAND2X1TS U2519 ( .A(n2051), .B(addWeight_16__add_biasesStored[1]), .Y(n161)
         );
  NAND2X1TS U2520 ( .A(n2051), .B(addWeight_16__add_biasesStored[0]), .Y(n169)
         );
  CLKBUFX2TS U2521 ( .A(n2032), .Y(n2052) );
  NAND2X1TS U2522 ( .A(n2052), .B(addWeight_15__add_biasesStored[1]), .Y(n151)
         );
  NAND2X1TS U2523 ( .A(n2052), .B(addWeight_15__add_biasesStored[0]), .Y(n159)
         );
  NAND2X1TS U2524 ( .A(n2033), .B(addWeight_14__add_biasesStored[1]), .Y(n141)
         );
  NAND2X1TS U2525 ( .A(n2033), .B(addWeight_14__add_biasesStored[0]), .Y(n149)
         );
  NAND2X1TS U2526 ( .A(n2044), .B(addWeight_13__add_biasesStored[1]), .Y(n131)
         );
  NAND2X1TS U2527 ( .A(n2044), .B(addWeight_13__add_biasesStored[0]), .Y(n139)
         );
  NAND2X1TS U2528 ( .A(n2055), .B(addWeight_10__add_biasesStored[1]), .Y(n101)
         );
  NAND2X1TS U2529 ( .A(n2040), .B(addWeight_10__add_biasesStored[0]), .Y(n109)
         );
  NAND2X1TS U2530 ( .A(n2056), .B(addWeight_9__add_biasesStored[1]), .Y(n91)
         );
  NAND2X1TS U2531 ( .A(n2043), .B(addWeight_9__add_biasesStored[0]), .Y(n99)
         );
  CLKBUFX2TS U2532 ( .A(n2034), .Y(n2063) );
  NAND2X1TS U2533 ( .A(n2063), .B(addWeight_8__add_biasesStored[1]), .Y(n81)
         );
  CLKBUFX2TS U2534 ( .A(n2034), .Y(n2066) );
  NAND2X1TS U2535 ( .A(n2066), .B(addWeight_8__add_biasesStored[0]), .Y(n89)
         );
  NAND2X1TS U2536 ( .A(n2057), .B(addWeight_7__add_biasesStored[1]), .Y(n71)
         );
  NAND2X1TS U2537 ( .A(n2041), .B(addWeight_7__add_biasesStored[0]), .Y(n79)
         );
  NAND2X1TS U2538 ( .A(n2058), .B(addWeight_6__add_biasesStored[1]), .Y(n61)
         );
  CLKBUFX2TS U2539 ( .A(n2035), .Y(n2062) );
  NAND2X1TS U2540 ( .A(n2062), .B(addWeight_6__add_biasesStored[0]), .Y(n69)
         );
  NAND2X1TS U2541 ( .A(n2070), .B(addWeight_5__add_biasesStored[1]), .Y(n51)
         );
  NAND2X1TS U2542 ( .A(n2060), .B(addWeight_5__add_biasesStored[0]), .Y(n59)
         );
  NAND2X1TS U2543 ( .A(n2060), .B(addWeight_4__add_biasesStored[1]), .Y(n41)
         );
  NAND2X1TS U2544 ( .A(n2065), .B(addWeight_4__add_biasesStored[0]), .Y(n49)
         );
  NAND2X1TS U2545 ( .A(n2036), .B(addWeight_3__add_biasesStored[1]), .Y(n31)
         );
  NAND2X1TS U2546 ( .A(n2036), .B(addWeight_3__add_biasesStored[0]), .Y(n39)
         );
  NAND2X1TS U2547 ( .A(n2043), .B(addWeight_0__add_biasesStored[1]), .Y(n1) );
  NAND2X1TS U2548 ( .A(n2046), .B(addWeight_0__add_biasesStored[0]), .Y(n9) );
  NAND2X1TS U2549 ( .A(n2057), .B(addWeight_31__add_biasesStored[3]), .Y(n315)
         );
  NAND2X1TS U2550 ( .A(n2036), .B(addWeight_30__add_biasesStored[3]), .Y(n305)
         );
  NAND2X1TS U2551 ( .A(n2069), .B(addWeight_29__add_biasesStored[3]), .Y(n295)
         );
  NAND2X1TS U2552 ( .A(n2053), .B(addWeight_24__add_biasesStored[3]), .Y(n245)
         );
  NAND2X1TS U2553 ( .A(n2038), .B(addWeight_23__add_biasesStored[3]), .Y(n235)
         );
  NAND2X1TS U2554 ( .A(n2045), .B(addWeight_22__add_biasesStored[3]), .Y(n225)
         );
  NAND2X1TS U2555 ( .A(n2047), .B(addWeight_21__add_biasesStored[3]), .Y(n215)
         );
  NAND2X1TS U2556 ( .A(n2047), .B(addWeight_20__add_biasesStored[3]), .Y(n205)
         );
  NAND2X1TS U2557 ( .A(n2048), .B(addWeight_19__add_biasesStored[3]), .Y(n195)
         );
  NAND2X1TS U2558 ( .A(n2049), .B(addWeight_18__add_biasesStored[3]), .Y(n185)
         );
  NAND2X1TS U2559 ( .A(n2037), .B(addWeight_17__add_biasesStored[3]), .Y(n175)
         );
  NAND2X1TS U2560 ( .A(n2038), .B(addWeight_16__add_biasesStored[3]), .Y(n165)
         );
  NAND2X1TS U2561 ( .A(n2039), .B(addWeight_15__add_biasesStored[3]), .Y(n155)
         );
  NAND2X1TS U2562 ( .A(n2053), .B(addWeight_14__add_biasesStored[3]), .Y(n145)
         );
  NAND2X1TS U2563 ( .A(n2054), .B(addWeight_13__add_biasesStored[3]), .Y(n135)
         );
  NAND2X1TS U2564 ( .A(n2055), .B(addWeight_10__add_biasesStored[3]), .Y(n105)
         );
  NAND2X1TS U2565 ( .A(n2040), .B(addWeight_9__add_biasesStored[3]), .Y(n95)
         );
  NAND2X1TS U2566 ( .A(n2061), .B(addWeight_8__add_biasesStored[3]), .Y(n85)
         );
  NAND2X1TS U2567 ( .A(n2066), .B(addWeight_7__add_biasesStored[3]), .Y(n75)
         );
  NAND2X1TS U2568 ( .A(n2041), .B(addWeight_6__add_biasesStored[3]), .Y(n65)
         );
  NAND2X1TS U2569 ( .A(n2058), .B(addWeight_5__add_biasesStored[3]), .Y(n55)
         );
  NAND2X1TS U2570 ( .A(n2059), .B(addWeight_4__add_biasesStored[3]), .Y(n45)
         );
  NAND2X1TS U2571 ( .A(n2059), .B(addWeight_3__add_biasesStored[3]), .Y(n35)
         );
  NAND2X1TS U2572 ( .A(n2042), .B(addWeight_2__add_biasesStored[3]), .Y(n25)
         );
  NAND2X1TS U2573 ( .A(n2041), .B(addWeight_31__add_biasesStored[2]), .Y(n313)
         );
  NAND2X1TS U2574 ( .A(n2042), .B(addWeight_30__add_biasesStored[2]), .Y(n303)
         );
  NAND2X1TS U2575 ( .A(n2070), .B(addWeight_29__add_biasesStored[2]), .Y(n293)
         );
  NAND2X1TS U2576 ( .A(n2043), .B(addWeight_27__add_biasesStored[2]), .Y(n273)
         );
  NAND2X1TS U2577 ( .A(n2044), .B(addWeight_25__add_biasesStored[2]), .Y(n253)
         );
  NAND2X1TS U2578 ( .A(n2052), .B(addWeight_24__add_biasesStored[2]), .Y(n243)
         );
  NAND2X1TS U2579 ( .A(n2050), .B(addWeight_23__add_biasesStored[2]), .Y(n233)
         );
  NAND2X1TS U2580 ( .A(n2045), .B(addWeight_22__add_biasesStored[2]), .Y(n223)
         );
  NAND2X1TS U2581 ( .A(n2046), .B(addWeight_21__add_biasesStored[2]), .Y(n213)
         );
  NAND2X1TS U2582 ( .A(n2047), .B(addWeight_20__add_biasesStored[2]), .Y(n203)
         );
  NAND2X1TS U2583 ( .A(n2048), .B(addWeight_19__add_biasesStored[2]), .Y(n193)
         );
  NAND2X1TS U2584 ( .A(n2049), .B(addWeight_18__add_biasesStored[2]), .Y(n183)
         );
  NAND2X1TS U2585 ( .A(n2050), .B(addWeight_17__add_biasesStored[2]), .Y(n173)
         );
  NAND2X1TS U2586 ( .A(n2051), .B(addWeight_16__add_biasesStored[2]), .Y(n163)
         );
  NAND2X1TS U2587 ( .A(n2052), .B(addWeight_15__add_biasesStored[2]), .Y(n153)
         );
  NAND2X1TS U2588 ( .A(n2053), .B(addWeight_14__add_biasesStored[2]), .Y(n143)
         );
  NAND2X1TS U2589 ( .A(n2054), .B(addWeight_13__add_biasesStored[2]), .Y(n133)
         );
  NAND2X1TS U2590 ( .A(n2055), .B(addWeight_10__add_biasesStored[2]), .Y(n103)
         );
  NAND2X1TS U2591 ( .A(n2056), .B(addWeight_9__add_biasesStored[2]), .Y(n93)
         );
  NAND2X1TS U2592 ( .A(n2063), .B(addWeight_8__add_biasesStored[2]), .Y(n83)
         );
  NAND2X1TS U2593 ( .A(n2057), .B(addWeight_7__add_biasesStored[2]), .Y(n73)
         );
  NAND2X1TS U2594 ( .A(n2058), .B(addWeight_6__add_biasesStored[2]), .Y(n63)
         );
  NAND2X1TS U2595 ( .A(n2062), .B(addWeight_5__add_biasesStored[2]), .Y(n53)
         );
  NAND2X1TS U2596 ( .A(n2059), .B(addWeight_4__add_biasesStored[2]), .Y(n43)
         );
  NAND2X1TS U2597 ( .A(n2060), .B(addWeight_3__add_biasesStored[2]), .Y(n33)
         );
  NAND2X1TS U2598 ( .A(n2061), .B(addWeight_27__add_biasesStored[3]), .Y(n275)
         );
  NAND2X1TS U2599 ( .A(n2063), .B(addWeight_0__add_biasesStored[2]), .Y(n3) );
  NAND2X1TS U2600 ( .A(n2062), .B(addWeight_29__add_biasesStored[0]), .Y(n299)
         );
  NAND2X1TS U2601 ( .A(n2067), .B(addWeight_11__add_biasesStored[0]), .Y(n119)
         );
  NAND2X1TS U2602 ( .A(n2062), .B(addWeight_1__add_biasesStored[2]), .Y(n13)
         );
  NAND2X1TS U2603 ( .A(n2063), .B(addWeight_0__add_biasesStored[3]), .Y(n5) );
  NAND2X1TS U2604 ( .A(n2066), .B(addWeight_28__add_biasesStored[0]), .Y(n289)
         );
  CLKBUFX2TS U2605 ( .A(n2064), .Y(n2073) );
  NAND2X1TS U2606 ( .A(n2073), .B(addWeight_11__add_biasesStored[2]), .Y(n113)
         );
  NAND2X1TS U2607 ( .A(n2073), .B(addWeight_11__add_biasesStored[1]), .Y(n111)
         );
  NAND2X1TS U2608 ( .A(n2068), .B(addWeight_26__add_biasesStored[0]), .Y(n269)
         );
  NAND2X1TS U2609 ( .A(n2071), .B(addWeight_12__add_biasesStored[2]), .Y(n123)
         );
  NAND2X1TS U2610 ( .A(n2067), .B(addWeight_26__add_biasesStored[2]), .Y(n263)
         );
  NAND2X1TS U2611 ( .A(n2068), .B(addWeight_12__add_biasesStored[0]), .Y(n129)
         );
  NAND2X1TS U2612 ( .A(n2074), .B(addWeight_28__add_biasesStored[1]), .Y(n281)
         );
  NAND2X1TS U2613 ( .A(n2065), .B(addWeight_2__add_biasesStored[0]), .Y(n29)
         );
  NAND2X1TS U2614 ( .A(n2071), .B(addWeight_25__add_biasesStored[3]), .Y(n255)
         );
  NAND2X1TS U2615 ( .A(n2073), .B(addWeight_11__add_biasesStored[3]), .Y(n115)
         );
  NAND2X1TS U2616 ( .A(n2066), .B(addWeight_28__add_biasesStored[2]), .Y(n283)
         );
  NAND2X1TS U2617 ( .A(n2067), .B(addWeight_26__add_biasesStored[3]), .Y(n265)
         );
  NAND2X1TS U2618 ( .A(n2068), .B(addWeight_12__add_biasesStored[1]), .Y(n121)
         );
  NAND2X1TS U2619 ( .A(n2069), .B(addWeight_1__add_biasesStored[3]), .Y(n15)
         );
  NAND2X1TS U2620 ( .A(n2074), .B(addWeight_28__add_biasesStored[3]), .Y(n285)
         );
  NAND2X1TS U2621 ( .A(n2070), .B(addWeight_2__add_biasesStored[1]), .Y(n21)
         );
  NAND2X1TS U2622 ( .A(n2071), .B(addWeight_12__add_biasesStored[3]), .Y(n125)
         );
  NAND2X1TS U2623 ( .A(n2072), .B(addWeight_1__add_biasesStored[1]), .Y(n11)
         );
  NAND2X1TS U2624 ( .A(n2073), .B(addWeight_26__add_biasesStored[1]), .Y(n261)
         );
  NAND2X1TS U2625 ( .A(n2074), .B(addWeight_1__add_biasesStored[0]), .Y(n19)
         );
  CLKBUFX2TS U2626 ( .A(n2136), .Y(n2076) );
  CLKBUFX2TS U2627 ( .A(n2076), .Y(n2357) );
  CLKBUFX2TS U2628 ( .A(n2076), .Y(n2356) );
  CLKBUFX2TS U2629 ( .A(n2075), .Y(n2078) );
  CLKBUFX2TS U2630 ( .A(n2078), .Y(n2334) );
  CLKBUFX2TS U2631 ( .A(n2076), .Y(n2355) );
  CLKBUFX2TS U2632 ( .A(n2077), .Y(n2348) );
  CLKBUFX2TS U2633 ( .A(n2077), .Y(n2347) );
  CLKBUFX2TS U2634 ( .A(n2077), .Y(n2346) );
  CLKBUFX2TS U2635 ( .A(n2078), .Y(n2335) );
  CLKBUFX2TS U2636 ( .A(n2078), .Y(n2331) );
  CLKBUFX2TS U2637 ( .A(n2079), .Y(n2080) );
  CLKBUFX2TS U2638 ( .A(n2080), .Y(n2093) );
  NAND2BXLTS U2639 ( .AN(addWeight_30__add_biasesStored[1]), .B(n2093), .Y(
        n302) );
  CLKBUFX2TS U2640 ( .A(clr), .Y(n2083) );
  CLKBUFX2TS U2641 ( .A(n2083), .Y(n2084) );
  CLKBUFX2TS U2642 ( .A(n2084), .Y(n2107) );
  NAND2BXLTS U2643 ( .AN(addWeight_25__add_biasesStored[0]), .B(n2107), .Y(
        n260) );
  CLKBUFX2TS U2644 ( .A(n2079), .Y(n2091) );
  CLKBUFX2TS U2645 ( .A(n2091), .Y(n2116) );
  NAND2BXLTS U2646 ( .AN(addWeight_27__add_biasesStored[1]), .B(n2116), .Y(
        n272) );
  CLKBUFX2TS U2647 ( .A(n2079), .Y(n2086) );
  CLKBUFX2TS U2648 ( .A(n2086), .Y(n2119) );
  NAND2BXLTS U2649 ( .AN(addWeight_2__add_biasesStored[2]), .B(n2119), .Y(n24)
         );
  NAND2BXLTS U2650 ( .AN(addWeight_25__add_biasesStored[1]), .B(n2107), .Y(
        n252) );
  CLKBUFX2TS U2651 ( .A(n2083), .Y(n2085) );
  CLKBUFX2TS U2652 ( .A(n2085), .Y(n2106) );
  NAND2BXLTS U2653 ( .AN(addWeight_27__add_biasesStored[0]), .B(n2106), .Y(
        n280) );
  CLKBUFX2TS U2654 ( .A(n2085), .Y(n2110) );
  NAND2BXLTS U2655 ( .AN(addWeight_2__add_biasesStored[0]), .B(n2110), .Y(n30)
         );
  CLKBUFX2TS U2656 ( .A(n2084), .Y(n2111) );
  NAND2BXLTS U2657 ( .AN(addWeight_26__add_biasesStored[0]), .B(n2111), .Y(
        n270) );
  CLKBUFX2TS U2658 ( .A(n2080), .Y(n2117) );
  NAND2BXLTS U2659 ( .AN(addWeight_24__add_biasesStored[0]), .B(n2117), .Y(
        n250) );
  CLKBUFX2TS U2660 ( .A(n2080), .Y(n2092) );
  NAND2BXLTS U2661 ( .AN(addWeight_29__add_biasesStored[1]), .B(n2092), .Y(
        n292) );
  CLKBUFX2TS U2662 ( .A(n2084), .Y(n2105) );
  NAND2BXLTS U2663 ( .AN(addWeight_28__add_biasesStored[0]), .B(n2105), .Y(
        n290) );
  NAND2BXLTS U2664 ( .AN(addWeight_24__add_biasesStored[1]), .B(n2117), .Y(
        n242) );
  CLKBUFX2TS U2665 ( .A(n2081), .Y(n2088) );
  CLKBUFX2TS U2666 ( .A(n2088), .Y(n2099) );
  NAND2BXLTS U2667 ( .AN(addWeight_11__add_biasesStored[0]), .B(n2099), .Y(
        n120) );
  CLKBUFX2TS U2668 ( .A(n2080), .Y(n2102) );
  NAND2BXLTS U2669 ( .AN(addWeight_30__add_biasesStored[0]), .B(n2102), .Y(
        n310) );
  CLKBUFX2TS U2670 ( .A(n2081), .Y(n2096) );
  CLKBUFX2TS U2671 ( .A(n2096), .Y(n2104) );
  NAND2BXLTS U2672 ( .AN(addWeight_12__add_biasesStored[0]), .B(n2104), .Y(
        n130) );
  NAND2BXLTS U2673 ( .AN(addWeight_28__add_biasesStored[1]), .B(n2111), .Y(
        n282) );
  NAND2BXLTS U2674 ( .AN(addWeight_23__add_biasesStored[1]), .B(n2093), .Y(
        n232) );
  CLKBUFX2TS U2675 ( .A(n2091), .Y(n2125) );
  NAND2BXLTS U2676 ( .AN(addWeight_31__add_biasesStored[0]), .B(n2125), .Y(
        n320) );
  NAND2BXLTS U2677 ( .AN(addWeight_31__add_biasesStored[1]), .B(n2116), .Y(
        n312) );
  CLKBUFX2TS U2678 ( .A(n2085), .Y(n2115) );
  NAND2BXLTS U2679 ( .AN(addWeight_1__add_biasesStored[0]), .B(n2115), .Y(n20)
         );
  NAND2BXLTS U2680 ( .AN(addWeight_26__add_biasesStored[1]), .B(n2105), .Y(
        n262) );
  NAND2BXLTS U2681 ( .AN(addWeight_29__add_biasesStored[0]), .B(n2107), .Y(
        n300) );
  NAND2BXLTS U2682 ( .AN(addWeight_12__add_biasesStored[1]), .B(n2104), .Y(
        n122) );
  NAND2BXLTS U2683 ( .AN(addWeight_11__add_biasesStored[1]), .B(n2099), .Y(
        n112) );
  NAND2BXLTS U2684 ( .AN(addWeight_2__add_biasesStored[1]), .B(n2110), .Y(n22)
         );
  NAND2BXLTS U2685 ( .AN(addWeight_1__add_biasesStored[1]), .B(n2115), .Y(n12)
         );
  CLKBUFX2TS U2686 ( .A(n2091), .Y(n2101) );
  CLKBUFX2TS U2687 ( .A(n2086), .Y(n2094) );
  NAND2BXLTS U2688 ( .AN(addWeight_4__add_biasesStored[2]), .B(n2094), .Y(n44)
         );
  CLKBUFX2TS U2689 ( .A(n2086), .Y(n2127) );
  NAND2BXLTS U2690 ( .AN(addWeight_5__add_biasesStored[2]), .B(n2127), .Y(n54)
         );
  CLKBUFX2TS U2691 ( .A(n2082), .Y(n2087) );
  CLKBUFX2TS U2692 ( .A(n2087), .Y(n2131) );
  NAND2BXLTS U2693 ( .AN(addWeight_6__add_biasesStored[2]), .B(n2131), .Y(n64)
         );
  CLKBUFX2TS U2694 ( .A(n2087), .Y(n2130) );
  NAND2BXLTS U2695 ( .AN(addWeight_7__add_biasesStored[2]), .B(n2130), .Y(n74)
         );
  CLKBUFX2TS U2696 ( .A(n2087), .Y(n2097) );
  NAND2BXLTS U2697 ( .AN(addWeight_8__add_biasesStored[2]), .B(n2097), .Y(n84)
         );
  CLKBUFX2TS U2698 ( .A(n2088), .Y(n2132) );
  NAND2BXLTS U2699 ( .AN(addWeight_9__add_biasesStored[2]), .B(n2132), .Y(n94)
         );
  CLKBUFX2TS U2700 ( .A(n2088), .Y(n2109) );
  NAND2BXLTS U2701 ( .AN(addWeight_10__add_biasesStored[2]), .B(n2109), .Y(
        n104) );
  CLKBUFX2TS U2702 ( .A(n2096), .Y(n2120) );
  NAND2BXLTS U2703 ( .AN(addWeight_13__add_biasesStored[2]), .B(n2120), .Y(
        n134) );
  CLKBUFX2TS U2704 ( .A(n2096), .Y(n2128) );
  NAND2BXLTS U2705 ( .AN(addWeight_14__add_biasesStored[2]), .B(n2128), .Y(
        n144) );
  CLKBUFX2TS U2706 ( .A(n2083), .Y(n2089) );
  CLKBUFX2TS U2707 ( .A(n2089), .Y(n2098) );
  NAND2BXLTS U2708 ( .AN(addWeight_15__add_biasesStored[2]), .B(n2098), .Y(
        n154) );
  CLKBUFX2TS U2709 ( .A(n2089), .Y(n2123) );
  NAND2BXLTS U2710 ( .AN(addWeight_16__add_biasesStored[2]), .B(n2123), .Y(
        n164) );
  CLKBUFX2TS U2711 ( .A(n2089), .Y(n2121) );
  NAND2BXLTS U2712 ( .AN(addWeight_17__add_biasesStored[2]), .B(n2121), .Y(
        n174) );
  CLKBUFX2TS U2713 ( .A(n2083), .Y(n2090) );
  CLKBUFX2TS U2714 ( .A(n2090), .Y(n2114) );
  NAND2BXLTS U2715 ( .AN(addWeight_18__add_biasesStored[2]), .B(n2114), .Y(
        n184) );
  CLKBUFX2TS U2716 ( .A(n2090), .Y(n2100) );
  NAND2BXLTS U2717 ( .AN(addWeight_19__add_biasesStored[2]), .B(n2100), .Y(
        n194) );
  CLKBUFX2TS U2718 ( .A(n2090), .Y(n2124) );
  NAND2BXLTS U2719 ( .AN(addWeight_20__add_biasesStored[2]), .B(n2124), .Y(
        n204) );
  NAND2BXLTS U2720 ( .AN(addWeight_21__add_biasesStored[2]), .B(n2125), .Y(
        n214) );
  NAND2BXLTS U2721 ( .AN(addWeight_22__add_biasesStored[2]), .B(n2101), .Y(
        n224) );
  NAND2BXLTS U2722 ( .AN(addWeight_23__add_biasesStored[2]), .B(n2102), .Y(
        n234) );
  NAND2BXLTS U2723 ( .AN(addWeight_24__add_biasesStored[2]), .B(n2092), .Y(
        n244) );
  CLKBUFX2TS U2724 ( .A(n2084), .Y(n2095) );
  NAND2BXLTS U2725 ( .AN(addWeight_25__add_biasesStored[2]), .B(n2095), .Y(
        n254) );
  CLKBUFX2TS U2726 ( .A(n2085), .Y(n2103) );
  NAND2BXLTS U2727 ( .AN(addWeight_27__add_biasesStored[2]), .B(n2103), .Y(
        n274) );
  NAND2BXLTS U2728 ( .AN(addWeight_29__add_biasesStored[2]), .B(n2092), .Y(
        n294) );
  NAND2BXLTS U2729 ( .AN(addWeight_30__add_biasesStored[2]), .B(n2093), .Y(
        n304) );
  NAND2BXLTS U2730 ( .AN(addWeight_31__add_biasesStored[2]), .B(n2116), .Y(
        n314) );
  NAND2BXLTS U2731 ( .AN(addWeight_2__add_biasesStored[3]), .B(n2119), .Y(n26)
         );
  CLKBUFX2TS U2732 ( .A(n2086), .Y(n2113) );
  NAND2BXLTS U2733 ( .AN(addWeight_3__add_biasesStored[3]), .B(n2113), .Y(n36)
         );
  NAND2BXLTS U2734 ( .AN(addWeight_4__add_biasesStored[3]), .B(n2094), .Y(n46)
         );
  CLKBUFX2TS U2735 ( .A(n2087), .Y(n2122) );
  NAND2BXLTS U2736 ( .AN(addWeight_5__add_biasesStored[3]), .B(n2122), .Y(n56)
         );
  NAND2BXLTS U2737 ( .AN(addWeight_6__add_biasesStored[3]), .B(n2131), .Y(n66)
         );
  NAND2BXLTS U2738 ( .AN(addWeight_7__add_biasesStored[3]), .B(n2130), .Y(n76)
         );
  NAND2BXLTS U2739 ( .AN(addWeight_8__add_biasesStored[3]), .B(n2097), .Y(n86)
         );
  CLKBUFX2TS U2740 ( .A(n2088), .Y(n2112) );
  NAND2BXLTS U2741 ( .AN(addWeight_9__add_biasesStored[3]), .B(n2112), .Y(n96)
         );
  NAND2BXLTS U2742 ( .AN(addWeight_10__add_biasesStored[3]), .B(n2109), .Y(
        n106) );
  NAND2BXLTS U2743 ( .AN(addWeight_13__add_biasesStored[3]), .B(n2120), .Y(
        n136) );
  NAND2BXLTS U2744 ( .AN(addWeight_14__add_biasesStored[3]), .B(n2128), .Y(
        n146) );
  NAND2BXLTS U2745 ( .AN(addWeight_15__add_biasesStored[3]), .B(n2098), .Y(
        n156) );
  CLKBUFX2TS U2746 ( .A(n2089), .Y(n2129) );
  NAND2BXLTS U2747 ( .AN(addWeight_16__add_biasesStored[3]), .B(n2129), .Y(
        n166) );
  NAND2BXLTS U2748 ( .AN(addWeight_17__add_biasesStored[3]), .B(n2121), .Y(
        n176) );
  NAND2BXLTS U2749 ( .AN(addWeight_18__add_biasesStored[3]), .B(n2114), .Y(
        n186) );
  NAND2BXLTS U2750 ( .AN(addWeight_28__add_biasesStored[7]), .B(n2095), .Y(
        n288) );
  NAND2BXLTS U2751 ( .AN(addWeight_19__add_biasesStored[3]), .B(n2100), .Y(
        n196) );
  CLKBUFX2TS U2752 ( .A(n2090), .Y(n2126) );
  NAND2BXLTS U2753 ( .AN(addWeight_20__add_biasesStored[3]), .B(n2126), .Y(
        n206) );
  CLKBUFX2TS U2754 ( .A(n2091), .Y(n2108) );
  NAND2BXLTS U2755 ( .AN(addWeight_21__add_biasesStored[3]), .B(n2108), .Y(
        n216) );
  NAND2BXLTS U2756 ( .AN(addWeight_22__add_biasesStored[3]), .B(n2108), .Y(
        n226) );
  NAND2BXLTS U2757 ( .AN(addWeight_3__add_biasesStored[2]), .B(n2113), .Y(n34)
         );
  NAND2BXLTS U2758 ( .AN(addWeight_23__add_biasesStored[3]), .B(n2102), .Y(
        n236) );
  NAND2BXLTS U2759 ( .AN(addWeight_24__add_biasesStored[3]), .B(n2092), .Y(
        n246) );
  NAND2BXLTS U2760 ( .AN(addWeight_28__add_biasesStored[3]), .B(n2095), .Y(
        n286) );
  NAND2BXLTS U2761 ( .AN(addWeight_29__add_biasesStored[3]), .B(n2117), .Y(
        n296) );
  NAND2BXLTS U2762 ( .AN(addWeight_30__add_biasesStored[3]), .B(n2108), .Y(
        n306) );
  NAND2BXLTS U2763 ( .AN(addWeight_31__add_biasesStored[3]), .B(n2125), .Y(
        n316) );
  NAND2BXLTS U2764 ( .AN(addWeight_27__add_biasesStored[3]), .B(n2106), .Y(
        n276) );
  NAND2BXLTS U2765 ( .AN(addWeight_0__add_biasesStored[0]), .B(n2093), .Y(n10)
         );
  NAND2BXLTS U2766 ( .AN(addWeight_0__add_biasesStored[1]), .B(n2109), .Y(n2)
         );
  NAND2BXLTS U2767 ( .AN(addWeight_3__add_biasesStored[0]), .B(n2119), .Y(n40)
         );
  NAND2BXLTS U2768 ( .AN(addWeight_26__add_biasesStored[3]), .B(n2106), .Y(
        n266) );
  NAND2BXLTS U2769 ( .AN(addWeight_3__add_biasesStored[1]), .B(n2113), .Y(n32)
         );
  NAND2BXLTS U2770 ( .AN(addWeight_4__add_biasesStored[0]), .B(n2094), .Y(n50)
         );
  NAND2BXLTS U2771 ( .AN(addWeight_4__add_biasesStored[1]), .B(n2094), .Y(n42)
         );
  NAND2BXLTS U2772 ( .AN(addWeight_25__add_biasesStored[3]), .B(n2095), .Y(
        n256) );
  NAND2BXLTS U2773 ( .AN(addWeight_5__add_biasesStored[0]), .B(n2127), .Y(n60)
         );
  NAND2BXLTS U2774 ( .AN(addWeight_5__add_biasesStored[1]), .B(n2127), .Y(n52)
         );
  NAND2BXLTS U2775 ( .AN(addWeight_6__add_biasesStored[0]), .B(n2122), .Y(n70)
         );
  CLKBUFX2TS U2776 ( .A(n2096), .Y(n2118) );
  NAND2BXLTS U2777 ( .AN(addWeight_12__add_biasesStored[3]), .B(n2118), .Y(
        n126) );
  NAND2BXLTS U2778 ( .AN(addWeight_6__add_biasesStored[1]), .B(n2122), .Y(n62)
         );
  NAND2BXLTS U2779 ( .AN(addWeight_7__add_biasesStored[0]), .B(n2131), .Y(n80)
         );
  NAND2BXLTS U2780 ( .AN(addWeight_7__add_biasesStored[1]), .B(n2130), .Y(n72)
         );
  NAND2BXLTS U2781 ( .AN(addWeight_11__add_biasesStored[3]), .B(n2099), .Y(
        n116) );
  NAND2BXLTS U2782 ( .AN(addWeight_8__add_biasesStored[0]), .B(n2097), .Y(n90)
         );
  NAND2BXLTS U2783 ( .AN(addWeight_8__add_biasesStored[1]), .B(n2097), .Y(n82)
         );
  NAND2BXLTS U2784 ( .AN(addWeight_9__add_biasesStored[0]), .B(n2132), .Y(n100) );
  NAND2BXLTS U2785 ( .AN(addWeight_1__add_biasesStored[3]), .B(n2110), .Y(n16)
         );
  NAND2BXLTS U2786 ( .AN(addWeight_9__add_biasesStored[1]), .B(n2132), .Y(n92)
         );
  NAND2BXLTS U2787 ( .AN(addWeight_10__add_biasesStored[0]), .B(n2112), .Y(
        n110) );
  NAND2BXLTS U2788 ( .AN(addWeight_10__add_biasesStored[1]), .B(n2112), .Y(
        n102) );
  NAND2BXLTS U2789 ( .AN(addWeight_0__add_biasesStored[3]), .B(n2103), .Y(n6)
         );
  NAND2BXLTS U2790 ( .AN(addWeight_13__add_biasesStored[0]), .B(n2118), .Y(
        n140) );
  NAND2BXLTS U2791 ( .AN(addWeight_13__add_biasesStored[1]), .B(n2118), .Y(
        n132) );
  NAND2BXLTS U2792 ( .AN(addWeight_14__add_biasesStored[0]), .B(n2120), .Y(
        n150) );
  NAND2BXLTS U2793 ( .AN(addWeight_28__add_biasesStored[2]), .B(n2111), .Y(
        n284) );
  NAND2BXLTS U2794 ( .AN(addWeight_14__add_biasesStored[1]), .B(n2128), .Y(
        n142) );
  NAND2BXLTS U2795 ( .AN(addWeight_15__add_biasesStored[0]), .B(n2098), .Y(
        n160) );
  NAND2BXLTS U2796 ( .AN(addWeight_15__add_biasesStored[1]), .B(n2098), .Y(
        n152) );
  NAND2BXLTS U2797 ( .AN(addWeight_26__add_biasesStored[2]), .B(n2105), .Y(
        n264) );
  NAND2BXLTS U2798 ( .AN(addWeight_16__add_biasesStored[0]), .B(n2123), .Y(
        n170) );
  NAND2BXLTS U2799 ( .AN(addWeight_16__add_biasesStored[1]), .B(n2123), .Y(
        n162) );
  NAND2BXLTS U2800 ( .AN(addWeight_17__add_biasesStored[0]), .B(n2129), .Y(
        n180) );
  NAND2BXLTS U2801 ( .AN(addWeight_12__add_biasesStored[2]), .B(n2104), .Y(
        n124) );
  NAND2BXLTS U2802 ( .AN(addWeight_17__add_biasesStored[1]), .B(n2129), .Y(
        n172) );
  NAND2BXLTS U2803 ( .AN(addWeight_18__add_biasesStored[0]), .B(n2121), .Y(
        n190) );
  NAND2BXLTS U2804 ( .AN(addWeight_18__add_biasesStored[1]), .B(n2114), .Y(
        n182) );
  NAND2BXLTS U2805 ( .AN(addWeight_11__add_biasesStored[2]), .B(n2099), .Y(
        n114) );
  NAND2BXLTS U2806 ( .AN(addWeight_19__add_biasesStored[0]), .B(n2100), .Y(
        n200) );
  NAND2BXLTS U2807 ( .AN(addWeight_19__add_biasesStored[1]), .B(n2100), .Y(
        n192) );
  NAND2BXLTS U2808 ( .AN(addWeight_20__add_biasesStored[0]), .B(n2124), .Y(
        n210) );
  NAND2BXLTS U2809 ( .AN(addWeight_1__add_biasesStored[2]), .B(n2115), .Y(n14)
         );
  NAND2BXLTS U2810 ( .AN(addWeight_20__add_biasesStored[1]), .B(n2124), .Y(
        n202) );
  NAND2BXLTS U2811 ( .AN(addWeight_21__add_biasesStored[0]), .B(n2126), .Y(
        n220) );
  NAND2BXLTS U2812 ( .AN(addWeight_21__add_biasesStored[1]), .B(n2126), .Y(
        n212) );
  NAND2BXLTS U2813 ( .AN(addWeight_0__add_biasesStored[2]), .B(n2103), .Y(n4)
         );
  NAND2BXLTS U2814 ( .AN(addWeight_22__add_biasesStored[0]), .B(n2101), .Y(
        n230) );
  NAND2BXLTS U2815 ( .AN(addWeight_22__add_biasesStored[1]), .B(n2101), .Y(
        n222) );
  NAND2BXLTS U2816 ( .AN(addWeight_23__add_biasesStored[7]), .B(n2102), .Y(
        n238) );
  NAND2BXLTS U2817 ( .AN(addWeight_31__add_biasesStored[7]), .B(n2103), .Y(
        n318) );
  NAND2BXLTS U2818 ( .AN(addWeight_11__add_biasesStored[7]), .B(n2104), .Y(
        n118) );
  NAND2BXLTS U2819 ( .AN(addWeight_27__add_biasesStored[7]), .B(n2105), .Y(
        n278) );
  NAND2BXLTS U2820 ( .AN(addWeight_26__add_biasesStored[7]), .B(n2106), .Y(
        n268) );
  NAND2BXLTS U2821 ( .AN(addWeight_24__add_biasesStored[7]), .B(n2107), .Y(
        n248) );
  NAND2BXLTS U2822 ( .AN(addWeight_22__add_biasesStored[7]), .B(n2108), .Y(
        n228) );
  NAND2BXLTS U2823 ( .AN(addWeight_10__add_biasesStored[7]), .B(n2109), .Y(
        n108) );
  NAND2BXLTS U2824 ( .AN(addWeight_1__add_biasesStored[7]), .B(n2110), .Y(n18)
         );
  NAND2BXLTS U2825 ( .AN(addWeight_25__add_biasesStored[7]), .B(n2111), .Y(
        n258) );
  NAND2BXLTS U2826 ( .AN(addWeight_9__add_biasesStored[7]), .B(n2112), .Y(n98)
         );
  NAND2BXLTS U2827 ( .AN(addWeight_3__add_biasesStored[7]), .B(n2113), .Y(n38)
         );
  NAND2BXLTS U2828 ( .AN(addWeight_18__add_biasesStored[7]), .B(n2114), .Y(
        n188) );
  NAND2BXLTS U2829 ( .AN(addWeight_0__add_biasesStored[7]), .B(n2115), .Y(n8)
         );
  NAND2BXLTS U2830 ( .AN(addWeight_21__add_biasesStored[7]), .B(n2116), .Y(
        n218) );
  NAND2BXLTS U2831 ( .AN(addWeight_29__add_biasesStored[7]), .B(n2117), .Y(
        n298) );
  NAND2BXLTS U2832 ( .AN(addWeight_12__add_biasesStored[7]), .B(n2118), .Y(
        n128) );
  NAND2BXLTS U2833 ( .AN(addWeight_2__add_biasesStored[7]), .B(n2119), .Y(n28)
         );
  NAND2BXLTS U2834 ( .AN(addWeight_13__add_biasesStored[7]), .B(n2120), .Y(
        n138) );
  NAND2BXLTS U2835 ( .AN(addWeight_17__add_biasesStored[7]), .B(n2121), .Y(
        n178) );
  NAND2BXLTS U2836 ( .AN(addWeight_5__add_biasesStored[7]), .B(n2122), .Y(n58)
         );
  NAND2BXLTS U2837 ( .AN(addWeight_15__add_biasesStored[7]), .B(n2123), .Y(
        n158) );
  NAND2BXLTS U2838 ( .AN(addWeight_19__add_biasesStored[7]), .B(n2124), .Y(
        n198) );
  NAND2BXLTS U2839 ( .AN(addWeight_30__add_biasesStored[7]), .B(n2125), .Y(
        n308) );
  NAND2BXLTS U2840 ( .AN(addWeight_20__add_biasesStored[7]), .B(n2126), .Y(
        n208) );
  NAND2BXLTS U2841 ( .AN(addWeight_4__add_biasesStored[7]), .B(n2127), .Y(n48)
         );
  NAND2BXLTS U2842 ( .AN(addWeight_14__add_biasesStored[7]), .B(n2128), .Y(
        n148) );
  NAND2BXLTS U2843 ( .AN(addWeight_16__add_biasesStored[7]), .B(n2129), .Y(
        n168) );
  NAND2BXLTS U2844 ( .AN(addWeight_7__add_biasesStored[7]), .B(n2130), .Y(n78)
         );
  NAND2BXLTS U2845 ( .AN(addWeight_6__add_biasesStored[7]), .B(n2131), .Y(n68)
         );
  NAND2BXLTS U2846 ( .AN(addWeight_8__add_biasesStored[7]), .B(n2132), .Y(n88)
         );
  CLKBUFX2TS U2847 ( .A(n2134), .Y(n2360) );
  CLKBUFX2TS U2848 ( .A(n2299), .Y(n2133) );
  CLKBUFX2TS U2849 ( .A(n2133), .Y(n2364) );
  CLKBUFX2TS U2850 ( .A(n2133), .Y(n2365) );
  CLKBUFX2TS U2851 ( .A(n2133), .Y(n2366) );
  CLKBUFX2TS U2852 ( .A(n2134), .Y(n2349) );
  CLKBUFX2TS U2853 ( .A(n2135), .Y(n2342) );
  CLKBUFX2TS U2854 ( .A(n2135), .Y(n2340) );
  AOI2BB1X1TS U2855 ( .A0N(n2385), .A1N(n2138), .B0(n2137), .Y(
        addWeight_24__add_s[0]) );
  AOI2BB1X1TS U2856 ( .A0N(sumOut[152]), .A1N(n2140), .B0(n2139), .Y(
        addWeight_19__add_s[0]) );
  AOI2BB1X1TS U2857 ( .A0N(sumOut[80]), .A1N(n2142), .B0(n2141), .Y(
        addWeight_10__add_s[0]) );
  AOI2BB1X1TS U2858 ( .A0N(sumOut[184]), .A1N(n2144), .B0(n2143), .Y(
        addWeight_23__add_s[0]) );
  AOI2BB1X1TS U2859 ( .A0N(sumOut[200]), .A1N(n2146), .B0(n2145), .Y(
        addWeight_25__add_s[0]) );
  AOI2BB1X1TS U2860 ( .A0N(sumOut[176]), .A1N(n2148), .B0(n2147), .Y(
        addWeight_22__add_s[0]) );
  AOI2BB1X1TS U2861 ( .A0N(sumOut[168]), .A1N(n2150), .B0(n2149), .Y(
        addWeight_21__add_s[0]) );
  AOI2BB1X1TS U2862 ( .A0N(sumOut[216]), .A1N(n366), .B0(n2151), .Y(
        addWeight_27__add_s[0]) );
  AOI2BB1X1TS U2863 ( .A0N(sumOut[0]), .A1N(n2153), .B0(n2152), .Y(
        addWeight_0__add_s[0]) );
  AOI2BB1X1TS U2864 ( .A0N(n2394), .A1N(n2155), .B0(n2154), .Y(
        addWeight_20__add_s[0]) );
  AOI2BB1X1TS U2865 ( .A0N(sumOut[240]), .A1N(n2157), .B0(n2156), .Y(
        addWeight_30__add_s[0]) );
  AOI2BB1X1TS U2866 ( .A0N(sumOut[16]), .A1N(n2159), .B0(n2158), .Y(
        addWeight_2__add_s[0]) );
  AOI2BB1X1TS U2867 ( .A0N(sumOut[208]), .A1N(n2161), .B0(n2160), .Y(
        addWeight_26__add_s[0]) );
  AOI2BB1X1TS U2868 ( .A0N(sumOut[224]), .A1N(n2164), .B0(n2163), .Y(
        addWeight_28__add_s[0]) );
  AOI2BB1X1TS U2869 ( .A0N(sumOut[232]), .A1N(n2172), .B0(n2171), .Y(
        addWeight_29__add_s[0]) );
  INVX2TS U2870 ( .A(n2173), .Y(n2175) );
  NAND2X1TS U2871 ( .A(n2175), .B(n2174), .Y(n2176) );
  XNOR2X1TS U2872 ( .A(n2177), .B(n2176), .Y(addWeight_3__add_s[2]) );
  INVX2TS U2873 ( .A(n2178), .Y(n2180) );
  NAND2X1TS U2874 ( .A(n2180), .B(n2179), .Y(n2181) );
  XNOR2X1TS U2875 ( .A(n2182), .B(n2181), .Y(addWeight_4__add_s[2]) );
  INVX2TS U2876 ( .A(n2183), .Y(n2185) );
  NAND2X1TS U2877 ( .A(n2185), .B(n2184), .Y(n2186) );
  XNOR2X1TS U2878 ( .A(n2187), .B(n2186), .Y(addWeight_5__add_s[2]) );
  INVX2TS U2879 ( .A(n2188), .Y(n2190) );
  NAND2X1TS U2880 ( .A(n2190), .B(n2189), .Y(n2191) );
  XNOR2X1TS U2881 ( .A(n2192), .B(n2191), .Y(addWeight_6__add_s[2]) );
  INVX2TS U2882 ( .A(n2193), .Y(n2195) );
  NAND2X1TS U2883 ( .A(n2195), .B(n2194), .Y(n2196) );
  XNOR2X1TS U2884 ( .A(n2197), .B(n2196), .Y(addWeight_7__add_s[2]) );
  INVX2TS U2885 ( .A(n2198), .Y(n2200) );
  NAND2X1TS U2886 ( .A(n2200), .B(n2199), .Y(n2201) );
  XNOR2X1TS U2887 ( .A(n2202), .B(n2201), .Y(addWeight_8__add_s[2]) );
  INVX2TS U2888 ( .A(n2203), .Y(n2205) );
  NAND2X1TS U2889 ( .A(n2205), .B(n2204), .Y(n2206) );
  XNOR2X1TS U2890 ( .A(n2207), .B(n2206), .Y(addWeight_9__add_s[2]) );
  INVX2TS U2891 ( .A(n2208), .Y(n2210) );
  NAND2X1TS U2892 ( .A(n2210), .B(n2209), .Y(n2211) );
  XNOR2X1TS U2893 ( .A(n2212), .B(n2211), .Y(addWeight_10__add_s[2]) );
  INVX2TS U2894 ( .A(n2213), .Y(n2215) );
  NAND2X1TS U2895 ( .A(n2215), .B(n2214), .Y(n2216) );
  XNOR2X1TS U2896 ( .A(n2217), .B(n2216), .Y(addWeight_13__add_s[2]) );
  INVX2TS U2897 ( .A(n2218), .Y(n2220) );
  NAND2X1TS U2898 ( .A(n2220), .B(n2219), .Y(n2221) );
  XNOR2X1TS U2899 ( .A(n2222), .B(n2221), .Y(addWeight_14__add_s[2]) );
  INVX2TS U2900 ( .A(n2223), .Y(n2225) );
  NAND2X1TS U2901 ( .A(n2225), .B(n2224), .Y(n2226) );
  XNOR2X1TS U2902 ( .A(n2227), .B(n2226), .Y(addWeight_15__add_s[2]) );
  INVX2TS U2903 ( .A(n2228), .Y(n2230) );
  NAND2X1TS U2904 ( .A(n2230), .B(n2229), .Y(n2231) );
  XNOR2X1TS U2905 ( .A(n2232), .B(n2231), .Y(addWeight_16__add_s[2]) );
  INVX2TS U2906 ( .A(n2233), .Y(n2235) );
  XNOR2X1TS U2907 ( .A(n2236), .B(n2237), .Y(addWeight_25__add_s[2]) );
  INVX2TS U2908 ( .A(n2238), .Y(n2240) );
  NAND2X1TS U2909 ( .A(n2240), .B(n2239), .Y(n2241) );
  XNOR2X1TS U2910 ( .A(n2242), .B(n2241), .Y(addWeight_24__add_s[2]) );
  INVX2TS U2911 ( .A(n2243), .Y(n2245) );
  NAND2X1TS U2912 ( .A(n2245), .B(n2244), .Y(n2246) );
  XNOR2X1TS U2913 ( .A(n2247), .B(n2246), .Y(addWeight_20__add_s[2]) );
  INVX2TS U2914 ( .A(n2248), .Y(n2250) );
  NAND2X1TS U2915 ( .A(n2250), .B(n2249), .Y(n2251) );
  XNOR2X1TS U2916 ( .A(n2252), .B(n2251), .Y(addWeight_18__add_s[2]) );
  INVX2TS U2917 ( .A(n2253), .Y(n2255) );
  NAND2X1TS U2918 ( .A(n2255), .B(n2254), .Y(n2256) );
  XNOR2X1TS U2919 ( .A(n2257), .B(n2256), .Y(addWeight_31__add_s[2]) );
  INVX2TS U2920 ( .A(n2258), .Y(n2260) );
  NAND2X1TS U2921 ( .A(n2260), .B(n2259), .Y(n2261) );
  XNOR2X1TS U2922 ( .A(n2262), .B(n2261), .Y(addWeight_30__add_s[2]) );
  INVX2TS U2923 ( .A(n2263), .Y(n2265) );
  NAND2X1TS U2924 ( .A(n2265), .B(n2264), .Y(n2266) );
  XNOR2X1TS U2925 ( .A(n2267), .B(n2266), .Y(addWeight_27__add_s[2]) );
  INVX2TS U2926 ( .A(n2268), .Y(n2270) );
  NAND2X1TS U2927 ( .A(n2270), .B(n2269), .Y(n2271) );
  XNOR2X1TS U2928 ( .A(n2272), .B(n2271), .Y(addWeight_17__add_s[2]) );
  INVX2TS U2929 ( .A(n2273), .Y(n2275) );
  NAND2X1TS U2930 ( .A(n2275), .B(n2274), .Y(n2276) );
  XNOR2X1TS U2931 ( .A(n2277), .B(n2276), .Y(addWeight_23__add_s[2]) );
  INVX2TS U2932 ( .A(n2278), .Y(n2280) );
  NAND2X1TS U2933 ( .A(n2280), .B(n2279), .Y(n2281) );
  XNOR2X1TS U2934 ( .A(n2282), .B(n2281), .Y(addWeight_21__add_s[2]) );
  INVX2TS U2935 ( .A(n2283), .Y(n2285) );
  NAND2X1TS U2936 ( .A(n2285), .B(n2284), .Y(n2286) );
  XNOR2X1TS U2937 ( .A(n2287), .B(n2286), .Y(addWeight_19__add_s[2]) );
  INVX2TS U2938 ( .A(n2288), .Y(n2290) );
  NAND2X1TS U2939 ( .A(n2290), .B(n2289), .Y(n2291) );
  XNOR2X1TS U2940 ( .A(n2292), .B(n2291), .Y(addWeight_22__add_s[2]) );
  INVX2TS U2941 ( .A(n462), .Y(n2295) );
  NAND2X1TS U2942 ( .A(n2295), .B(n2294), .Y(n2296) );
  XNOR2X1TS U2943 ( .A(n2297), .B(n2296), .Y(addWeight_2__add_s[2]) );
endmodule

