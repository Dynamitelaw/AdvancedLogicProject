`include "EntireNetwork.v"


module Generated_TestBench ;
	//Instantiate modules
	reg reset = 0;
	reg clk;
	reg inputsInbound = 0;
	reg predictionRecieved = 0;
	reg inputPixel;
	reg weightWriteEnable;
	reg biasWriteEnable;
	reg LayerWriteSelect;
	reg [9:0] WriteAddressSelect;
	reg [`WRITE_IN_BIT_WIDTH-1:0] writeIn;
	
	wire predictionReady;
	wire readyForInputs;
	wire [3:0] predictionOut;
	NN_Controler controller(
		//Inputs
	 	.reset(reset), 
	 	.masterClk(clk), 
	 	.inputsInbound(inputsInbound), 
	 	.predictionRecieved(predictionRecieved),
	 	.inputPixel(inputPixel), 
	 	.weightWriteEnable(weightWriteEnable), 
	 	.biasWriteEnable(biasWriteEnable), 
	 	.LayerWriteSelect(LayerWriteSelect), 
	 	.WriteAddressSelect(WriteAddressSelect), 
	 	.writeIn(writeIn),
		//Outputs
	 	.predictionReady(predictionReady), 
	 	.readyForInputs(readyForInputs),
	 	.predictionOut(predictionOut)
	);
	
	reg[783:0] inputVectors [19:0];  //InputVectors
	reg currentInputIndex = 0;

	initial
	begin
		clk = 0;
		#1

		//=================================
		//--Load in weights and Biases--
		//=================================

		//Layer 1 Weights
		#1
		LayerWriteSelect = 0;
		#1
		#2
		WriteAddressSelect <= 10'b0;  //node 0
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_00000_00001_00001_00001_00000_00001_00000_11111_00000_00001_11111_00000_00001_00001_00000_00001_00001_11111_00001_00001_00000_11111_11110_00000_00010_00001_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1;  //node 1
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00001_11110_00000_11111_11111_00010_00000_00000_00001_00000_00000_00001_11111_11111_00000_11110_00001_00001_11111_00000_00001_00001_11111_00000_11111_11111_00001_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b10;  //node 2
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_11111_11111_00000_11111_00000_00000_00000_11111_00001_00001_00000_00010_11111_00001_00000_11111_00001_11110_11111_00001_00000_00001_00000_11111_11111_11111_11111_11111;

		#2
		WriteAddressSelect <= 10'b11;  //node 3
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00001_00000_11110_00001_11111_00001_11111_00000_00000_00000_11111_00000_00000_00000_00001_11111_11111_11111_00000_00001_11101_00001_00000_00000_11111_11111_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b100;  //node 4
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00001_00000_00000_11111_00001_00000_11111_00010_11111_11111_00001_00001_00010_11110_00010_00001_11110_00001_11111_11110_00000_00000_00000_00010_11110_00001_00000_00001_00000_11110;

		#2
		WriteAddressSelect <= 10'b101;  //node 5
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00001_00000_11111_00000_00000_11111_00000_00000_00000_00000_11111_00010_00001_00000_11111_11111_00001_00001_00010_00000_00010_00010_11111_11111_00000_11111_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b110;  //node 6
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00001_00000_11110_00010_00010_00010_00010_11111_00001_00000_00001_11111_00001_00001_00000_11111_00001_00000_00001_00000_11110_00000_11111_00000_11111_00000_00000_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b111;  //node 7
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00000_11111_11110_00001_11111_11110_00000_00001_00000_00000_00001_11111_00001_11111_00000_00000_11111_00000_11111_00010_00000_00000_00010_00001_11111_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b1000;  //node 8
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_00000_00000_00000_11111_00001_00001_00001_11111_00001_00001_00000_00001_00000_11111_00000_00001_11111_00001_00001_11111_00001_11110_00001_00001_00000_00000_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1001;  //node 9
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_00000_00001_11111_00000_00000_00000_00000_00001_00000_11111_00010_00001_11110_11111_11111_00000_00010_00000_11110_00001_00001_11110_00001_00000_00001_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010;  //node 10
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_00000_00000_00000_11111_00001_11111_00000_11111_11111_11110_00001_00000_11101_00010_00000_00001_11111_00001_00000_00000_00000_00001_11111_00001_00000_11111_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b1011;  //node 11
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00010_11111_11111_11111_11111_00000_11111_11111_00000_11111_00010_00000_00000_00001_00001_11111_11110_00001_00001_00010_00001_00000_11111_11111_11111_00010_00001_00000_11110;

		#2
		WriteAddressSelect <= 10'b1100;  //node 12
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11111_00001_11111_11111_00000_00000_11111_00010_11110_00001_00000_00000_00000_11110_11111_11110_00000_00001_00001_11111_00010_11111_11111_00001_00000_00000_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1101;  //node 13
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00010_00001_11111_00000_11111_00000_00000_00000_00001_00000_11110_00000_11111_00000_11110_00001_00000_00000_11111_11111_00001_00000_00001_11111_00001_00001_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1110;  //node 14
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_00001_00001_00001_00000_11111_00000_11111_00000_00001_00010_11111_00010_00000_11110_00000_00000_00000_11111_00010_00000_00000_00000_00010_00000_11111_11111_11111_11110_00000;

		#2
		WriteAddressSelect <= 10'b1111;  //node 15
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00001_00001_00001_11111_00000_11111_00000_00010_00000_11110_00001_00000_00001_11111_00001_00001_00000_00000_11111_00001_00000_00000_00001_00001_00010_00000_00010_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b10000;  //node 16
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11111_00001_00000_11110_00000_00000_00001_00001_00000_00001_11110_11111_00001_00001_00010_11111_00001_00000_00000_00010_00000_00001_00000_00000_11111_11110_11110_00001_00001;

		#2
		WriteAddressSelect <= 10'b10001;  //node 17
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_11111_00000_00000_11111_00000_11110_11111_00000_00000_00000_00001_11110_11111_11111_00000_11111_00010_00010_11111_11111_00001_11111_00000_00010_00001_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b10010;  //node 18
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00000_00001_11111_00010_11111_00001_00000_00000_00000_00001_11111_11111_11111_00001_00001_00010_00001_00000_11111_00000_00010_11111_00000_11111_00010_11111_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b10011;  //node 19
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00010_00000_11111_00000_11111_11111_11111_11110_11111_11110_00000_00001_00000_11111_11111_11111_00000_00000_00000_00000_00000_00001_11110_11111_11111_11111_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b10100;  //node 20
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_00010_00001_00001_00000_11110_11111_00000_11110_00001_11111_11111_00001_11111_00001_00000_00001_11110_00000_00000_00000_00001_00000_11111_00000_11111_00000_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b10101;  //node 21
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11111_00000_00000_00001_00010_00000_00000_00010_00000_00001_00000_11111_00001_00000_00010_11110_00000_11111_00001_00001_00000_00000_11111_00001_00001_00000_11110_00000_11111;

		#2
		WriteAddressSelect <= 10'b10110;  //node 22
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00001_00000_00010_00000_00000_00000_00001_11110_00001_00000_00000_11111_11110_00001_00001_00000_00000_00001_11111_00001_11111_00000_00001_00000_00010_11111_11110_00010_00001;

		#2
		WriteAddressSelect <= 10'b10111;  //node 23
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00000_11111_00001_00000_00001_11111_00000_00001_00000_00010_11111_00000_00001_00010_11111_00000_00000_00000_00000_11111_00001_00001_00001_00010_00001_11110_00010_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b11000;  //node 24
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00010_00001_00000_11110_11111_00000_00010_11111_11111_00000_00000_00001_00001_00000_11111_11111_11111_11111_11111_00000_00000_00001_00000_00000_11111_00001_00001_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b11001;  //node 25
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_00000_11111_00000_11111_00000_11111_00000_00001_00000_11111_00000_00001_00000_00000_11110_11110_00000_00000_00000_00001_11110_00001_11111_00000_00000_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b11010;  //node 26
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_00000_00000_11111_00000_11111_00001_00001_11111_00000_00000_11111_11111_00000_00000_11111_00000_11111_11111_00010_00001_00000_00000_00001_00000_11111_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b11011;  //node 27
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00001_11110_00001_11111_00001_00001_11111_00001_00000_00000_00001_00000_00001_00010_00001_11111_00010_00000_00000_00000_00000_11111_00000_11111_00000_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b11100;  //node 28
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00000_11111_00001_00001_00001_11111_11110_11111_00001_00001_00000_00001_00000_11111_11111_11111_00000_00001_11111_00001_00000_00000_00001_11111_11111_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b11101;  //node 29
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00001_11111_00000_00000_00001_00010_00001_00001_11111_00001_00000_00000_00000_11111_11111_00010_00000_11111_00001_00000_00000_11111_00000_00000_00001_11111_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b11110;  //node 30
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_00001_11111_00001_00000_11111_00001_00000_00001_00000_11111_11111_00000_00010_11111_00010_00000_11111_00000_00000_11111_11110_00001_00001_11110_00000_00000_11110_00000_00000;

		#2
		WriteAddressSelect <= 10'b11111;  //node 31
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_00001_11111_11111_11111_00000_11110_00001_00001_11111_00001_11111_11111_00010_00001_11111_00000_00000_00000_00001_11111_00000_00010_11111_00000_00000_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b100000;  //node 32
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00010_00001_00000_11111_00000_11111_00000_00000_00001_00010_00001_11111_11111_00000_11111_11111_11111_11111_00000_11111_00000_00000_00010_11111_00000_00000_00010_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b100001;  //node 33
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_11111_00001_11111_00000_00001_00000_00000_00000_00000_11111_00001_00001_00001_00000_11111_00001_00001_00000_00010_00000_00001_00000_00001_00000_00000_00000_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b100010;  //node 34
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_11110_00000_00000_11110_00000_11111_00000_11111_00000_00000_11111_00000_00000_00001_00001_00010_00001_11111_00010_00000_11110_11110_00001_11110_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b100011;  //node 35
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_11111_00000_00000_11111_00000_00000_00000_00000_11111_11111_00001_11111_00000_11111_11111_11111_11111_00000_00001_00000_00010_00010_00000_00000_11111_00001_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b100100;  //node 36
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00001_00000_00000_00001_00001_00000_00000_00000_00000_00001_00001_11111_00001_00000_11110_00010_00000_00010_11111_00000_11111_00000_00000_11111_00001_00001_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b100101;  //node 37
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_11110_00010_11111_11110_00001_00000_11111_00000_11111_00000_00001_00000_00001_00000_00001_11111_11110_00001_00000_11111_00000_00010_00000_00000_11111_11111_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b100110;  //node 38
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_00000_11111_00000_00001_11111_00000_00000_00001_00001_11111_00001_00000_00000_00000_00001_00000_11111_00001_11110_11110_00000_00000_11111_00000_00000_11111_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b100111;  //node 39
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_11111_00001_00000_11111_00000_00000_11111_00001_11111_00001_11111_00000_00000_00010_00001_00000_00000_00000_00000_00000_00000_11111_00001_11111_00000_00000_00001_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b101000;  //node 40
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00010_11111_11111_00000_11111_00001_11111_00000_00010_11111_00001_00000_00000_00001_00000_00000_00000_00000_11110_00010_00000_00010_11111_11110_00000_00000_11110_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b101001;  //node 41
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00010_11111_00001_00000_11111_00000_11111_00000_00000_00000_00000_00000_11110_00000_00010_11111_00000_00000_00000_00000_00001_00000_00000_00010_11111_11111_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b101010;  //node 42
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_00001_00000_00001_11111_11111_00001_00001_00000_00000_11111_00001_11111_00001_00000_00010_00000_11111_11110_00010_00000_00000_00001_00000_00001_11111_00010_11110_00000_00000_00010;

		#2
		WriteAddressSelect <= 10'b101011;  //node 43
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00000_00010_00001_00001_00001_00000_11111_00000_00000_00000_00000_00000_00001_11111_00000_00000_11111_11111_11111_00001_00000_00001_11111_11111_00010_00001_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b101100;  //node 44
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00010_11111_11110_00001_11111_00010_11111_00000_00000_00000_00000_11111_00000_00000_00001_11111_00001_11110_00001_00000_00001_00000_00000_00000_11111_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b101101;  //node 45
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00001_11111_11110_00001_00000_00001_11111_00000_00000_11111_00000_00001_00001_00001_11111_00000_00000_00000_00001_00000_11111_00001_00000_00001_11111_00001_00000_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b101110;  //node 46
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00000_00001_00001_00000_00001_11110_00000_11111_00001_11111_00000_00001_00001_11111_11111_11111_00001_11111_00000_00000_00000_11111_00010_00000_11111_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b101111;  //node 47
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11111_00000_00001_00000_00000_00000_00001_00000_00001_00000_11111_00001_00000_11111_00000_11111_00001_00001_00000_00000_00000_00001_00000_00000_11111_00010_00000_11110_00001;

		#2
		WriteAddressSelect <= 10'b110000;  //node 48
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_11111_00001_00010_11111_11111_11110_11110_00000_00000_11111_11111_11111_00001_00000_11110_00000_00010_00000_11111_00000_11111_00001_00000_00000_00000_00000_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b110001;  //node 49
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_11110_00001_00001_00000_00001_00000_00001_11110_11111_00001_00000_00001_00000_00000_00000_00000_11111_11111_00000_11111_11111_00000_00000_00000_00000_00000_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b110010;  //node 50
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00001_11110_00001_00001_11111_00000_00000_11111_00000_11111_11111_00001_11110_00001_11111_11111_00001_00000_00000_00010_00000_00010_00000_00001_00000_11110_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b110011;  //node 51
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_00000_11111_00000_11111_00001_11111_11111_00001_11111_00001_00001_11110_00001_00001_00010_00001_00010_00000_00000_00001_11111_11111_00010_00010_00000_00000_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b110100;  //node 52
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11111_00001_00010_11111_11110_00010_00000_00001_00000_11111_11111_00000_00001_00001_11111_00001_11111_11111_00000_00000_00000_00000_00001_00001_00001_11111_11111_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b110101;  //node 53
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_11111_00001_11111_00000_11111_00000_00000_00001_00000_00000_11111_11111_11111_00000_00001_00001_11111_00001_00000_11111_00000_11111_00000_11111_00000_00000_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b110110;  //node 54
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_11111_00001_00000_00001_11111_11111_11110_00001_11111_11111_00000_00000_00001_00000_00001_00000_11111_00001_11111_00000_00001_11111_11110_11111_00000_11111_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b110111;  //node 55
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_11111_00000_00001_11111_00000_11111_00000_11111_00001_00000_00001_11111_00001_11110_00001_00001_00000_00001_00001_00001_11111_00000_00000_11111_00000_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b111000;  //node 56
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_00001_11111_11111_00000_00001_00000_11111_00001_00001_00000_00000_00010_00001_00010_00000_00001_00001_00001_11110_11111_00000_11110_11110_00001_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b111001;  //node 57
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00001_00000_00000_00000_00001_00000_00000_00001_11110_00000_00000_00000_00000_00010_00001_00000_00001_00001_00000_11111_11111_11111_11111_11111_11111_00000_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b111010;  //node 58
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_00000_00001_00001_00000_00001_00000_00000_00001_00001_00000_00000_00000_00000_00000_11110_00000_00000_11110_00000_00000_11111_00001_00000_00000_11111_00000_00010_11111_00010;

		#2
		WriteAddressSelect <= 10'b111011;  //node 59
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00001_00001_11111_00000_11111_00000_00001_00000_00000_00000_00001_00000_11111_00000_11111_11110_00010_00000_00000_00001_11111_11111_00000_00000_11110_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b111100;  //node 60
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00001_00000_11111_11111_11111_00000_11111_11111_11111_11111_00001_00000_00010_11111_00000_00001_11111_11110_00000_00001_00000_00000_11110_00000_00010_00001_11110_00001_00001;

		#2
		WriteAddressSelect <= 10'b111101;  //node 61
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00010_00000_00000_00001_11110_00000_00001_00000_11111_00000_00001_00001_00000_11111_00000_00001_11110_00001_11111_00000_00001_11111_00001_11110_00000_00000_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b111110;  //node 62
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_11111_00001_00001_11111_00000_11111_00001_00000_00000_11110_00000_00000_11110_00000_00001_11111_00010_00001_11111_00000_00000_11111_00001_00000_00000_00001_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b111111;  //node 63
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00001_11111_00001_00000_00000_00001_11111_11111_00000_00000_00001_00001_11111_00000_11110_00001_00000_00000_00000_11110_00001_11111_00000_00000_11111_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1000000;  //node 64
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_00000_00001_00001_00000_00001_00000_00001_00000_00001_11111_00000_00001_00001_11111_00000_11111_11111_00010_00001_11110_00001_00001_11111_00001_11111_11111_11110_00000;

		#2
		WriteAddressSelect <= 10'b1000001;  //node 65
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_00010_00000_11110_00001_11111_00001_11111_00001_11110_00001_00001_00001_00000_00000_00001_11111_00001_00001_00001_00000_00000_11111_11111_11110_00000_00001_00000_11110_11110;

		#2
		WriteAddressSelect <= 10'b1000010;  //node 66
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00000_11111_00000_00000_11111_00001_00010_11111_00000_00001_00001_00001_11110_00000_00000_00001_00001_00001_11110_11111_00010_11110_11111_11111_00000_00001_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1000011;  //node 67
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_00010_00000_00000_11110_00001_00000_00001_00000_00000_00010_00001_00001_11111_00001_00001_00001_00000_11111_00001_11110_00000_00001_00000_00000_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b1000100;  //node 68
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00000_00001_00001_00000_00001_00001_11110_11111_00000_00000_11111_00001_00000_00000_00001_00001_00010_00000_00000_00001_11111_00000_00000_00001_00000_11111_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1000101;  //node 69
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00000_11111_00000_00000_11111_00000_00001_00010_00000_11111_11111_00000_00000_00000_00000_00000_00000_00001_00001_00000_00001_00000_00000_11111_11111_00001_11111_00010_00001_00010;

		#2
		WriteAddressSelect <= 10'b1000110;  //node 70
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00010_00000_11111_11111_00000_11111_11111_00000_00000_00000_00000_00000_00000_00010_00000_00000_00000_00001_00001_00000_11111_11111_00000_00000_00000_11111_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b1000111;  //node 71
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_11111_00000_11111_00001_11110_11111_00000_00001_00000_11110_00001_11111_11111_00001_00001_00000_11110_00001_11111_00000_00000_00000_00000_11111_00000_11110_11111_11110;

		#2
		WriteAddressSelect <= 10'b1001000;  //node 72
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_00001_00001_00000_00001_00000_00001_00000_11111_00000_00000_00000_00000_11111_00001_11110_00000_11111_00001_00000_11111_00001_11111_00000_00000_00001_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b1001001;  //node 73
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_11111_00000_11111_00000_11111_00001_00000_00000_00000_00000_00000_11111_00000_00000_00000_11110_11111_00000_00001_11110_00010_11111_00000_11111_11110_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001010;  //node 74
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_00010_00001_00001_00000_00000_00001_00001_00000_00010_11111_00000_11111_00000_00000_11111_11111_00001_00000_00001_00001_11110_11110_00000_11111_11111_11111_11111_00010_00010;

		#2
		WriteAddressSelect <= 10'b1001011;  //node 75
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_00001_11110_00001_00000_11110_11111_00010_00000_00010_11111_00000_00001_11111_00001_00000_00000_00001_00000_00000_11111_00000_11110_11111_00001_00000_11110_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b1001100;  //node 76
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_00010_00010_00001_00001_00001_00000_00000_11111_11110_00001_00000_00001_11111_00001_00000_00001_00001_11111_11110_11111_00000_11111_00000_00000_00000_00001_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b1001101;  //node 77
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00001_00000_00010_11110_00000_00001_00000_11111_00000_11111_00001_11111_00000_00000_00001_11111_00001_00001_00000_00000_11111_00001_00000_00010_00000_11111_00000_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001110;  //node 78
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00010_11111_00001_00000_00000_00000_00000_00000_00000_00001_11111_11111_00000_11111_11111_11111_00001_00000_00000_00001_00000_11111_00000_00000_11110_00000_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001111;  //node 79
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11101_00010_00000_11111_00001_00000_00001_00001_11111_00000_00000_11111_00000_00001_00001_00000_00001_00000_11110_11111_00000_00000_11111_00000_00000_00000_00001_00000_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b1010000;  //node 80
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_11111_00000_00000_00001_00001_00000_00000_00000_11111_00001_11111_00001_11111_00000_00000_11111_11110_11111_00001_00000_11111_00001_11111_11111_00001_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1010001;  //node 81
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_00000_00000_11111_11111_00000_00001_11111_11110_11111_00001_00000_00000_00000_00000_00000_00001_11111_00010_00000_00000_00001_00001_00001_00010_00000_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1010010;  //node 82
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_11111_11110_11111_00000_11111_11111_00001_00001_11111_00000_00001_00000_00001_00001_11111_00000_11111_00000_11111_00000_00000_00001_11111_00000_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010011;  //node 83
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_11110_11110_00000_00000_11111_00000_00000_00010_00001_00000_00000_00000_00000_11111_00000_00000_00000_11110_11111_00001_00001_00010_00010_11111_00001_00001_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010100;  //node 84
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_00000_11111_11111_00000_00000_11111_11110_11110_00010_00001_00000_11111_00001_00000_00000_00000_00000_00001_00000_00001_00000_11111_00001_00001_00000_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b1010101;  //node 85
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11111_11111_11111_00010_00000_00001_11110_00001_00000_00000_00000_00001_11110_11111_00000_00001_00000_11111_00000_00001_00000_00000_11110_11111_11111_00000_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1010110;  //node 86
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_11111_00000_00000_11111_00000_00001_00001_00001_11111_11111_11111_11111_00000_00001_00001_00000_00000_11110_00000_00000_00010_00000_00001_11111_00000_00000_11111_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b1010111;  //node 87
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_11111_00000_11111_11111_00001_00010_11111_00000_00001_11111_00000_00010_00001_11111_00001_00000_00000_00001_11111_11111_00000_00000_00000_00010_00001_11111_11110_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011000;  //node 88
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00001_00001_00000_11111_00000_00000_00001_00001_00001_00000_11111_00000_11111_11111_00001_11111_11110_00000_00000_00010_11111_00000_00010_00000_00001_00001_11111_11111_11111;

		#2
		WriteAddressSelect <= 10'b1011001;  //node 89
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11110_00001_11110_00000_00001_00000_00010_11110_00000_00000_11110_00001_11111_00000_00000_00010_00010_11110_00000_00000_00000_00001_11111_00000_00000_11111_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011010;  //node 90
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_00001_00000_11111_00000_00000_00001_00000_00000_00000_00000_11101_00010_11110_00000_00001_00001_00000_00000_00001_00001_00000_00010_00001_00000_00000_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1011011;  //node 91
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00001_00000_00000_00000_11110_00000_00001_11110_00010_00010_11111_00000_00000_11110_00000_00000_11111_00001_00010_00000_00001_00001_00001_00001_11110_00000_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011100;  //node 92
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_11110_00000_00000_00000_00001_11110_00000_00001_00000_11111_00001_11111_00000_00001_11111_11110_11111_00001_00001_11111_00001_11111_00000_00001_00000_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011101;  //node 93
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00010_00001_11111_00001_00001_00000_11111_00000_11110_00010_00000_00000_00000_11111_00001_00000_00000_00000_00010_00001_00001_11111_00000_11111_11111_00001_00000_00010_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011110;  //node 94
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_11110_00001_00000_00001_00000_11111_11111_00001_00001_11111_00000_11111_00000_11111_11110_11111_00000_00000_11111_00000_00001_00000_00001_00000_11111_00000_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011111;  //node 95
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00001_00000_00000_00001_00001_00001_00001_00001_00000_00001_00001_11111_00000_11111_00001_00001_00000_00000_00001_00001_00000_00001_00000_00000_00000_00001_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1100000;  //node 96
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11111_11111_00010_00001_11111_00001_11111_00000_00000_00000_11110_11110_00000_11111_00001_00000_11111_00001_11111_00010_00001_11111_11111_11111_00010_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1100001;  //node 97
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00010_11110_11111_11111_11111_11111_00001_11111_11111_00001_00001_00000_11111_00001_00000_00001_11111_00000_00000_00000_00000_11111_11111_11111_00001_00000_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1100010;  //node 98
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_11111_00001_00000_00000_00000_11111_11110_00010_00000_00000_11110_00010_11110_00000_00000_11111_00000_11110_11111_11111_00000_11110_00010_00001_00001_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1100011;  //node 99
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00001_00000_00000_00001_00010_00000_00000_11110_11111_00000_00000_00001_00000_11111_11111_11110_00001_00001_00000_00001_00000_00001_00000_00000_00001_00001_00010_11111_11111;

		#2
		WriteAddressSelect <= 10'b1100100;  //node 100
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_11111_00000_11111_00000_11111_11111_00000_11111_11111_00010_00001_11110_00001_00000_11111_11110_00000_00001_00001_11111_00000_11111_11111_11111_00000_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1100101;  //node 101
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11110_11110_11111_00000_00001_11111_11111_00010_11111_00000_00010_00001_00000_00001_11111_00001_00001_00001_00001_00000_00000_00001_00000_00001_11110_00001_11111_00010_00000_00000;

		#2
		WriteAddressSelect <= 10'b1100110;  //node 102
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_00001_00000_00001_00010_11111_00000_00000_00000_11111_00000_00001_00001_11111_00000_00000_00000_00010_00001_00010_00000_00000_11110_00001_11111_00000_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b1100111;  //node 103
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_11111_11111_11110_00000_00001_00000_00000_11111_00000_00001_00000_00000_00001_00001_00000_00001_00000_11111_00000_11111_11111_00000_11111_00001_00001_11111_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1101000;  //node 104
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00001_00000_11110_00000_00000_00001_00001_00000_00001_00000_11111_00001_11110_00001_11111_00001_11110_00000_11111_00001_00001_11111_00001_11111_00001_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1101001;  //node 105
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_11111_11110_00000_00000_11111_00000_11111_00000_11111_11111_00000_00001_11111_00010_00001_00000_00000_00001_00001_00000_11111_00000_00000_00000_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1101010;  //node 106
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_00000_00000_00000_00010_11110_00010_11111_11110_11111_11110_11111_11111_00001_00001_11111_00010_00001_00001_00001_00001_00000_00001_11111_00001_00000_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1101011;  //node 107
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_00001_00000_00001_00000_00000_00001_00000_11111_00000_00000_00000_00000_11111_00000_00001_11110_00001_11111_00000_00000_00010_11111_00000_00001_00000_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1101100;  //node 108
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00001_00010_00000_11111_00000_00000_00001_11111_11111_00001_00001_00000_11111_00010_00000_00000_00010_11111_11110_00010_00001_00000_00000_11111_00001_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1101101;  //node 109
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_00001_00000_00000_00000_00001_00000_11111_00001_11111_11111_00010_11110_00001_00000_00000_00001_00000_11110_00001_00000_11111_00000_11111_00010_11111_11111_00001_00001_00010;

		#2
		WriteAddressSelect <= 10'b1101110;  //node 110
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_11110_00010_00000_00010_00001_11110_00001_00010_00000_11111_00000_11110_00001_00000_00001_11111_00000_11111_00001_00001_00001_00000_11111_00001_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1101111;  //node 111
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00010_11111_11111_00000_11111_11111_00000_00000_00000_00001_11111_00000_11111_00000_11111_11111_00000_00001_00000_00001_00000_00000_00000_00001_00000_00000_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1110000;  //node 112
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00001_11111_00000_11110_00000_11111_00000_00000_00000_00000_00000_00000_00000_11111_11111_11111_11111_11110_00001_00010_00000_00001_00000_00000_11110_00000_11111_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1110001;  //node 113
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_00001_11110_00001_00000_00000_00000_00001_11111_00000_11111_00001_00000_00000_00000_11111_00001_00000_00001_00000_11111_11111_11111_00000_11111_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b1110010;  //node 114
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00001_11111_00001_11111_00001_11111_11111_00010_11110_11111_00000_00000_00001_11111_00000_00000_00001_00010_00000_00010_00000_00001_11110_11110_00001_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1110011;  //node 115
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_00000_11111_11111_11110_00000_00001_00000_00000_11111_00000_11111_11111_11111_11111_00000_00000_11111_00010_00000_11111_00000_00000_00001_00000_00000_11110_00001_00010_00001;

		#2
		WriteAddressSelect <= 10'b1110100;  //node 116
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00010_00001_11111_11111_00010_00001_00001_11111_00000_00001_11111_11111_00000_00001_00001_00000_00000_11111_00001_00001_00000_11111_00010_00000_00000_00010_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1110101;  //node 117
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_00000_00001_00000_00001_00010_00000_11110_00000_00000_11111_00000_00000_00001_11111_00000_00000_00000_11110_00000_00001_11111_00001_11111_00000_00001_00000_11111_00000_11110;

		#2
		WriteAddressSelect <= 10'b1110110;  //node 118
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00001_00000_11111_11111_11111_00000_00000_11111_00010_00000_00001_11111_11111_00001_00001_00000_11111_00001_00000_11111_00001_00001_00000_00000_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1110111;  //node 119
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_00001_00000_00001_11110_00000_11111_00001_00000_00000_11111_00000_00001_00000_00001_11111_11110_11111_00000_00000_11110_00010_11111_11111_11111_11111_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1111000;  //node 120
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00010_11111_00001_00000_00010_00000_11111_00000_00000_00001_00000_00001_11111_00001_11110_00000_00000_11111_00001_11111_11111_00000_00000_11111_00000_00001_00000_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b1111001;  //node 121
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00000_00001_00001_00001_00000_11111_00000_00010_00010_11111_00000_11111_00000_11111_11111_11111_11111_00000_00001_00000_00001_00001_00000_00001_00000_00001_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b1111010;  //node 122
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_11111_00000_11111_00000_00001_11110_00000_11111_00001_00000_11111_00001_11111_00001_00001_00000_11111_11111_11111_00000_00001_11110_11111_11111_00001_00000_00000_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b1111011;  //node 123
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00010_11111_00010_00001_00000_00001_00000_00000_00001_11111_00000_00001_11111_00000_11111_00001_00001_00001_00001_11111_11111_11111_11110_00000_11110_00000_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1111100;  //node 124
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00001_00001_00000_00000_11111_11110_11110_11111_00000_00010_00000_11111_00001_00000_00000_11110_00000_00000_11110_00010_11111_11111_11111_00001_11111_00000_11111_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1111101;  //node 125
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11101_00000_00000_11110_00001_11111_00001_11111_00000_11111_00000_11111_11111_00000_11110_00001_11110_00001_00000_11110_11111_00010_00000_00000_00000_00010_00000_00001_00000_11111_11110;

		#2
		WriteAddressSelect <= 10'b1111110;  //node 126
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_00001_00000_00000_11111_00000_00001_00000_11111_00000_11111_11101_11111_00010_00001_11111_00000_00000_00000_00000_00001_11110_11111_11110_00000_11110_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1111111;  //node 127
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00010_00000_11111_00001_00000_00001_00000_00001_11111_11111_00001_00010_00000_11111_11110_11111_00001_00000_11111_11111_00000_00001_00001_00010_00000_00000_11111_00001_11110;

		#2
		WriteAddressSelect <= 10'b10000000;  //node 128
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_11111_00000_11111_11111_00000_11111_00000_11111_00000_00001_00000_00001_00000_11111_00000_00000_00001_00001_00000_00000_00000_11110_00001_00001_00000_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b10000001;  //node 129
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_11110_11110_00001_00001_00000_11111_11111_00001_00000_00000_11111_11111_11111_00000_00010_11111_00000_00000_00001_11110_11111_11111_00001_11110_11110_00001_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b10000010;  //node 130
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11110_00000_00010_11110_00001_00010_11111_00001_00000_00000_00010_00010_00010_00001_00001_00001_00010_00000_00001_11111_00010_00000_00000_00000_00000_11111_00000_11111_11111_11111;

		#2
		WriteAddressSelect <= 10'b10000011;  //node 131
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_11111_00000_00000_00000_00000_00001_11111_00000_00000_00001_00001_00000_11110_00010_00001_00000_00000_11110_11111_00000_00000_00000_11110_00000_00010_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b10000100;  //node 132
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11110_11111_00000_00000_00000_11110_11111_11111_00000_00000_00001_00001_00000_00001_00000_00000_00000_11111_11110_00001_00000_00001_11111_00001_11111_11111_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b10000101;  //node 133
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_00000_00000_00010_00000_11110_00001_00000_11111_00001_00010_00001_00010_00000_00000_11111_00000_11110_00010_00010_11111_00000_00001_00000_00000_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b10000110;  //node 134
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_00000_00000_00000_11111_00001_00000_00000_00000_11111_00010_00001_11111_00000_11111_00000_11111_00010_11111_00001_00001_00001_00001_00001_00001_00000_00001_00010;

		#2
		WriteAddressSelect <= 10'b10000111;  //node 135
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_11110_00000_00010_00000_11111_00000_00000_11111_00000_11111_00010_00000_11111_00000_00001_00010_00000_00000_11111_11111_11110_11111_11110_00000_11111_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b10001000;  //node 136
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00010_00001_00001_00000_11111_00000_11110_00000_00001_00001_00010_11110_11111_00000_00000_11111_11111_00000_11111_00001_00000_00001_00001_00000_00000_11111_00001_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b10001001;  //node 137
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11111_11110_11111_11111_11111_11111_00001_00001_11111_11110_00001_00001_00001_00010_00001_00010_00010_00010_00000_00001_00000_00000_00001_00001_11110_00000_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b10001010;  //node 138
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00001_11111_11110_00000_00001_11111_11110_00010_00000_00000_11111_00001_00001_00000_11111_00000_00000_11111_11111_00010_11110_00001_11111_00001_11111_11110_00001_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b10001011;  //node 139
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00001_11110_11111_00001_00010_00000_00001_11111_11111_00001_00000_00001_11111_00001_00010_00001_11111_00000_11110_00001_00000_00000_11111_00010_11111_00000_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b10001100;  //node 140
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00000_00000_00000_00001_00000_00000_00000_11111_00000_00000_11111_11111_00000_00001_00000_11111_00010_00000_00010_11111_00010_00000_00001_00000_00000_00000_00000_00000_11111_00010;

		#2
		WriteAddressSelect <= 10'b10001101;  //node 141
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_00001_11111_11111_00000_00000_11111_00001_00000_00000_11110_00000_00001_00001_00010_00001_11111_00000_00010_00010_00000_00001_00000_00000_00000_00001_11111_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b10001110;  //node 142
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00001_00001_00001_00000_00010_00001_11111_11111_00000_11111_00000_00001_00001_00000_00010_00000_00000_00000_00000_00000_00001_11110_11111_00010_00000_00001_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b10001111;  //node 143
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_11111_11111_11111_00001_11111_00010_00000_00001_00000_00000_00000_00000_00001_00000_00000_11111_00000_00000_00000_00000_00000_00000_11111_11111_11111_00001_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b10010000;  //node 144
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_11111_11110_11110_00000_00000_00001_00000_00000_00001_00001_00010_11111_11111_00001_00000_00010_11111_00000_00001_00001_00001_11110_00001_11111_00000_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b10010001;  //node 145
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_11111_00001_11111_00000_00001_00000_11111_11110_00001_00010_00000_00000_11111_00000_00000_11110_00000_00000_11111_11111_00001_00000_00000_00001_11111_00000_00000_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b10010010;  //node 146
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_11111_11111_00000_00000_00000_11111_00001_11111_00001_00001_11111_00000_00000_00000_00001_00000_00001_00010_11111_00001_11110_00001_00000_00000_00001_00000_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b10010011;  //node 147
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11111_00000_00001_00001_11111_11111_11111_11110_11110_00000_00000_00010_11110_00000_00000_00001_00000_11110_00001_00000_00000_00001_11111_00000_11111_00000_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b10010100;  //node 148
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00000_11110_00001_00000_00000_11111_00001_00000_00001_00000_00000_00000_00001_00000_11110_11111_00000_00000_00010_11110_00001_00001_11111_00000_00001_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b10010101;  //node 149
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11110_00010_00000_00001_11111_11111_00000_00000_00010_00001_00011_00001_11111_00010_00000_00000_00000_00000_00001_00000_11111_00001_11110_00000_00001_11111_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b10010110;  //node 150
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11110_00000_00001_11111_11111_11111_00000_11111_00000_00000_11111_11111_11111_00001_11111_11110_11111_00001_11111_11111_00000_00001_00001_11110_11110_00000_00000_00010_11111;

		#2
		WriteAddressSelect <= 10'b10010111;  //node 151
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11111_11111_00000_00001_11110_11110_00000_00000_00001_00001_00001_00001_11111_11110_00000_11101_00000_00010_00000_11111_00010_00000_00001_00000_00000_00000_00001_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b10011000;  //node 152
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11111_00000_00000_00000_11110_00000_11111_00001_00001_11111_11111_11101_11111_00001_11101_00000_00000_11111_11111_00000_11111_11111_00000_00000_11111_11111_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b10011001;  //node 153
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_11111_11111_00001_00001_00010_11111_00001_00001_00000_11111_11110_11110_00001_11100_00001_00001_11111_00000_00001_00010_00001_00000_00000_00001_00001_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b10011010;  //node 154
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11111_00000_00010_00000_00000_00010_00000_11110_00001_11101_11111_00000_11110_11111_11110_11110_11111_00000_00000_00000_00000_00000_00001_00000_00000_11111_00010_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b10011011;  //node 155
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_11111_11111_00001_11110_00000_11111_00001_00000_11111_11110_00001_00000_11111_00000_00000_00001_00000_11111_11110_11111_00000_00001_00001_00010_00001_00000_00000_00000_00001_00010;

		#2
		WriteAddressSelect <= 10'b10011100;  //node 156
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00000_00001_00001_00001_00000_11111_11111_11110_11110_11010_11110_11111_00000_00000_00010_11111_11111_00000_11111_00010_11110_00010_00000_11110_00000_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b10011101;  //node 157
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_00000_11111_11110_00000_00001_00001_11110_11110_11111_11110_11111_00000_00010_11110_00000_00000_11110_00001_11110_11110_00000_11110_00001_11111_11111_00010_11110_11111_00001;

		#2
		WriteAddressSelect <= 10'b10011110;  //node 158
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_11110_11110_00010_00000_00001_00010_00000_00001_11111_00001_00000_00001_00001_00001_11111_00001_00000_00001_00000_00000_11111_11110_00001_00001_11111_00000_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b10011111;  //node 159
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_00000_11111_00001_11110_00000_00001_00001_00000_00001_00000_00001_00001_00001_00000_11111_00001_00001_00001_00001_11111_00001_00000_11111_00000_00001_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b10100000;  //node 160
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00001_00001_00000_00001_11111_11111_00010_00000_11111_11110_11111_00001_00010_00000_00000_00001_11111_00001_11111_11111_00000_11111_11111_11110_00001_11110_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b10100001;  //node 161
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_00000_00000_00010_00000_00000_00000_00001_00001_11110_00001_00000_00001_00001_00001_00001_00000_00000_11111_00000_00000_11110_00000_00000_00000_00010_00010_11111_00000_11110;

		#2
		WriteAddressSelect <= 10'b10100010;  //node 162
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00001_00010_11111_00000_00001_11110_11111_00000_00001_00000_00001_11111_00001_00000_00001_00000_00000_00010_00000_00001_11110_00000_00010_00010_00001_00000_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b10100011;  //node 163
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11110_00001_11111_00000_11111_00001_00000_00000_00001_00010_00001_00001_00001_11111_11111_00001_00001_11111_00000_11110_00000_00000_00010_11111_11111_00001_00001_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b10100100;  //node 164
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_11111_00001_11111_00000_11110_11111_00000_00001_00001_11111_00000_00000_00001_00000_00000_00000_11111_00000_00010_00000_00000_11111_11111_00000_00000_00010_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b10100101;  //node 165
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00001_11111_00000_11111_11111_00000_11111_00010_00000_00001_00001_00000_00001_00001_00001_11111_11111_00001_00000_11110_00001_00000_00000_00000_11111_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b10100110;  //node 166
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00001_11111_11111_00000_00000_11111_11111_11111_00001_00010_00001_00000_00000_00000_00000_00001_00000_11111_00000_00001_11110_11110_00001_00001_11110_00000_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b10100111;  //node 167
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00000_00001_00000_00001_00000_11111_00010_00001_00000_00001_11111_00010_00000_00001_11111_00001_11111_00000_00000_00000_11111_11110_00001_11111_00000_00001_00001_11110_11111;

		#2
		WriteAddressSelect <= 10'b10101000;  //node 168
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_00001_11111_11111_00010_00001_00000_11111_00001_00001_00000_11111_00001_11111_00000_00010_00000_11111_11110_11111_00001_00001_00000_00001_00001_11111_00010_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b10101001;  //node 169
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_11111_00000_11111_00000_11111_11111_11111_00000_00001_11111_00000_00010_11110_11111_11111_11111_00001_11111_00010_00000_00000_00001_00001_00001_00001_00000_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b10101010;  //node 170
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_11110_00000_00000_11111_00001_11111_00001_00001_00001_00001_00000_11111_00000_00001_11111_00001_11111_00001_00000_00000_00000_00000_11111_00010_00000_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b10101011;  //node 171
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11110_00001_00010_00000_00000_11111_00000_00000_00000_00000_00000_00001_00000_11111_00000_00000_11111_00010_00000_00000_00000_11111_00000_11111_00000_00000_11110_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b10101100;  //node 172
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_00000_00000_00000_11111_11110_00001_00001_11110_00001_00001_11111_00010_11111_00001_00000_00000_11111_00000_00000_00000_00000_00001_11111_11111_00001_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b10101101;  //node 173
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11111_00001_11111_00000_00001_00000_00000_00000_11110_00001_00001_11111_00010_11111_11111_00001_00000_11111_00010_11111_11111_11111_00001_11111_00000_11110_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b10101110;  //node 174
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_00000_00000_00001_00000_00000_00010_00000_00001_00000_00000_00000_00001_11111_11111_00000_11111_11111_00000_00010_11111_00001_00001_00001_11110_00010_00001_11110_00001;

		#2
		WriteAddressSelect <= 10'b10101111;  //node 175
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_00001_00000_00001_00000_11110_00000_11111_00010_00000_11111_11111_00001_00000_11111_00001_11110_00000_11111_00001_00000_11110_00001_00001_00000_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b10110000;  //node 176
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00010_00001_11111_00000_11111_11110_00000_00000_00000_00001_11110_00001_00001_11111_00010_00000_00000_00010_00000_11111_11111_00000_00001_00001_11110_00001_00000_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b10110001;  //node 177
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00000_00000_00001_11110_00001_11111_11111_00010_00010_00000_00001_11111_00000_00000_00010_00001_11110_11111_00001_11111_00000_00010_00010_00000_11111_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b10110010;  //node 178
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_11111_11111_11111_11111_00001_11110_00000_00000_00011_11111_00000_00001_11111_00000_00000_00010_00000_11111_00001_11111_00000_11110_00001_11110_11111_00000_00010_00010_00001;

		#2
		WriteAddressSelect <= 10'b10110011;  //node 179
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00001_11111_00001_00000_11110_00000_00010_00000_00001_00010_11110_00010_00001_00000_00000_11110_11111_00001_00001_11111_00000_00000_00010_11111_11111_11111_11111_11111_00001_11110;

		#2
		WriteAddressSelect <= 10'b10110100;  //node 180
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11110_11111_00010_00000_11111_00000_00010_00000_00001_11111_00000_11110_11111_00000_11111_11100_11111_00000_11111_00000_11110_00010_11111_11110_11110_00001_00000_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b10110101;  //node 181
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_11110_00010_11111_00000_00000_00001_00000_00001_00001_11111_11111_11110_00001_00000_11011_00000_00000_11111_11111_00000_00000_00000_00010_11111_00000_00001_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b10110110;  //node 182
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_00010_11111_11110_00000_00000_00000_00001_11110_00000_11110_00010_11110_00000_11110_00000_00000_11111_00001_00001_11110_00000_00001_11110_00001_00000_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b10110111;  //node 183
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00001_00001_11111_11110_00001_00000_00000_11111_00000_00001_11110_11110_00001_00000_00001_00000_00000_00101_00001_11111_00000_00000_00001_11110_11111_00001_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b10111000;  //node 184
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_11111_00010_11110_11110_00010_00000_11101_11111_11110_00000_11110_11110_00001_00000_00001_11110_11111_00000_00000_00000_00001_00010_11111_00000_11111_00001_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b10111001;  //node 185
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11110_00001_00000_11110_11111_00001_00001_11110_11100_00000_00000_11111_00001_11111_11110_11111_11110_00000_11110_00000_11111_00010_00001_00000_00000_11111_00010_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b10111010;  //node 186
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11111_00001_11110_11111_00000_00000_11110_11111_11110_11111_00001_00011_11110_11111_00001_11111_11111_00010_00001_11110_00011_00001_00000_00000_11111_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b10111011;  //node 187
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00010_00000_11111_11110_00001_00000_00001_00001_00000_11110_00000_00010_00010_00010_11111_00000_11111_00001_00001_00000_11110_00001_11111_00000_00001_00000_00000_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b10111100;  //node 188
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00000_00000_11110_00010_00000_00001_00000_00000_11110_00000_00010_11111_00001_11111_11111_11111_00001_00010_00000_11101_00010_00010_00010_00000_11111_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b10111101;  //node 189
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_11111_11111_11111_11111_11111_00001_00001_00000_11111_11111_00001_00001_00010_00001_00000_00000_00010_11111_11110_11111_00000_00000_00001_00001_00011_00001_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b10111110;  //node 190
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00011_00000_00001_00001_00000_11111_00001_00010_11111_11111_00000_00010_00000_11111_00001_11111_11111_00000_00000_00000_11111_11111_00010_11110_11111_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b10111111;  //node 191
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00000_00000_11111_00000_00001_11110_00010_11111_00001_11111_00000_00001_00001_00000_00010_00001_00000_00010_11110_00010_11111_00000_00001_11111_11110_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b11000000;  //node 192
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00010_11110_00001_00001_00000_11111_00001_00000_00010_00001_00000_11111_11111_00000_00001_00000_11111_00000_11111_00001_11111_11111_00001_00000_00000_00000_11110_00000_11111;

		#2
		WriteAddressSelect <= 10'b11000001;  //node 193
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11110_00001_00000_00001_11111_00000_00000_00000_00001_11111_11111_00000_00001_11111_00000_00000_00001_00000_00001_11110_11111_11111_00000_11111_11110_00000_00010_00010_11111;

		#2
		WriteAddressSelect <= 10'b11000010;  //node 194
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00001_11111_11110_00000_00001_11110_11110_00000_11111_00000_00000_11110_11111_00000_00000_11111_11111_00000_00000_00001_00010_00000_00001_11111_00000_11111_00000_00010_11111_00001;

		#2
		WriteAddressSelect <= 10'b11000011;  //node 195
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00001_00000_00001_11111_00000_11110_00001_00000_00001_00010_00001_00000_11111_11111_11111_00000_00010_00000_00000_00001_11111_00000_00001_00001_11111_11110_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b11000100;  //node 196
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_00000_11111_00000_11111_00001_11111_11111_00000_11111_00000_11111_00000_11111_00001_00001_00010_00000_00000_00001_00000_00000_11111_11111_00000_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b11000101;  //node 197
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11111_11110_00000_11111_00001_00000_11110_00010_00000_00000_00000_00001_00000_11111_00000_11111_00000_00000_00000_00000_00000_00010_00000_11111_00000_00000_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b11000110;  //node 198
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00000_00000_00000_00000_00000_11111_11111_11111_00001_00000_11111_00001_00001_11111_00000_00010_00000_00001_00001_11111_00000_00001_00000_00001_00000_00001_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b11000111;  //node 199
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_11111_11110_11111_11111_11111_00001_00000_00000_00001_00010_00001_00000_00001_00001_00001_00001_00000_11111_00001_00000_00001_11111_00001_11111_11111_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b11001000;  //node 200
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11110_00000_00001_00001_00001_11111_00000_00000_00010_00000_11110_11111_00000_11111_11111_00000_11110_00000_00000_11110_00000_11111_00000_00000_00000_11111_11111_11110_11110;

		#2
		WriteAddressSelect <= 10'b11001001;  //node 201
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_00000_11111_00001_00010_00000_11110_00001_00001_00001_00000_00010_00001_00000_00010_00001_11111_11111_11111_00000_11110_11111_00010_00001_11111_00000_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b11001010;  //node 202
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_11111_11111_00000_00000_11111_11110_11111_00010_00001_00000_00001_00000_00001_00000_00001_11111_11111_00001_11111_00000_00001_00000_00000_00001_00001_11110_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b11001011;  //node 203
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_00000_00010_11111_00010_00000_00000_00001_00000_00001_11110_00010_11111_00000_00010_00001_11111_00000_00000_00000_11111_00000_11011_11110_00010_11111_11110_00010_11110_11110;

		#2
		WriteAddressSelect <= 10'b11001100;  //node 204
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00000_00001_00001_11110_00000_00000_00000_00000_11111_00000_11111_00000_00010_00001_11111_00001_00000_11111_00000_11111_00000_11111_00000_00001_00000_00011_00000_00001;

		#2
		WriteAddressSelect <= 10'b11001101;  //node 205
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00000_11111_00001_00001_11111_11111_00010_00001_00001_00001_11110_00001_00001_11111_00000_00001_00000_11111_00000_00000_00000_11111_11110_11111_00000_00000_00000_00010_11111_11111;

		#2
		WriteAddressSelect <= 10'b11001110;  //node 206
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_11110_11111_00000_00000_00001_00001_11111_00010_00010_11111_00001_00010_11111_00010_00000_00000_00010_11111_11110_00001_00000_00000_11111_11111_00000_00000_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b11001111;  //node 207
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00001_11111_11111_11111_00000_00010_00000_11111_00011_11111_00010_00000_00000_00001_11101_00000_00001_00000_11110_00001_00001_00010_00001_00000_11110_00001_00001_00001_00010;

		#2
		WriteAddressSelect <= 10'b11010000;  //node 208
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_11111_00000_00001_00001_00010_00010_11110_00001_00001_00001_11111_11110_00001_00010_11011_11111_00010_00000_00001_11111_11101_00000_00000_11110_00000_00001_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b11010001;  //node 209
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_00000_00010_11111_11111_00001_00010_00001_00010_00000_00000_11110_00001_11110_00000_11010_11111_00000_11111_00001_00010_00001_00000_00001_11111_00001_00001_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b11010010;  //node 210
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_11111_00000_00001_11111_00010_00001_00001_00010_11110_00001_11110_11110_00000_00001_11110_00000_11111_00001_11111_00000_00000_00001_00010_00010_00010_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b11010011;  //node 211
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_00000_00010_11101_11110_00010_00001_11111_00000_11110_00000_11111_11110_00001_00000_00010_00000_11111_00001_00001_11111_00000_11111_00000_11110_00000_00001_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b11010100;  //node 212
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_00000_00001_11111_11111_00010_00010_11100_00000_11111_11110_11110_11111_00001_11111_00010_00001_00000_00001_11111_00001_00000_00010_00010_11111_11111_11110_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b11010101;  //node 213
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11110_00000_00000_00001_00001_00010_11101_11110_00000_00000_11110_11111_00000_11111_11111_00000_11111_11111_00000_00000_00010_00001_00000_11111_00001_00010_00001_11110_11111;

		#2
		WriteAddressSelect <= 10'b11010110;  //node 214
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_00000_00001_11111_11111_00001_00001_11111_11101_11110_11110_00000_00000_11111_11111_11111_00000_11111_00000_00001_11111_00011_00010_00001_11110_11111_00001_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b11010111;  //node 215
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11111_11111_11111_00000_00000_11110_00001_00000_11110_00000_11110_00001_11110_11110_11110_00001_00000_00000_00001_00000_11110_00001_00000_00001_11111_11111_00000_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b11011000;  //node 216
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11111_00000_11111_00000_00000_11111_11111_00001_11111_11110_00000_00001_00001_00000_00001_11111_00001_00000_11110_11111_00001_00000_00001_00001_00000_00000_00010_00001_00000_11110;

		#2
		WriteAddressSelect <= 10'b11011001;  //node 217
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00001_11111_11111_00000_00000_00000_00010_00000_11110_00000_00001_00001_11111_11111_11111_11111_11111_00001_11111_00000_00000_00001_00000_11110_11111_00000_11110_00010_00000;

		#2
		WriteAddressSelect <= 10'b11011010;  //node 218
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00000_11111_00001_00001_11111_11111_00000_00000_11111_11111_00000_11111_00010_00000_00000_00000_00001_00000_11111_11111_11110_00001_00001_11111_00000_00001_00000_00000_00010;

		#2
		WriteAddressSelect <= 10'b11011011;  //node 219
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_11111_11111_00001_00000_00001_00000_11111_00001_00010_00010_11111_00000_00000_00010_00000_11111_00010_00001_00000_00001_11111_11110_00000_00000_00001_11111_11111_00000_00010;

		#2
		WriteAddressSelect <= 10'b11011100;  //node 220
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_11111_11111_00000_00000_00000_11111_00010_00001_00001_00001_11110_11110_00000_11111_11111_00010_11111_11111_00000_00010_00010_11111_11111_00000_00000_11111_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b11011101;  //node 221
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_11110_00000_00001_00001_00000_00001_11111_00001_11111_00001_00001_00000_00000_00000_00000_00010_00000_00001_00001_00001_00001_00000_00000_00001_00001_00001_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b11011110;  //node 222
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11111_00000_00000_00000_00000_00000_11111_00001_00010_00000_00000_00001_11111_00001_00000_00001_00000_00000_00000_00000_00000_11111_00001_11111_11111_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b11011111;  //node 223
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_11111_00000_00000_00000_00010_00000_11110_11111_11111_11111_00001_11110_00000_00001_00000_00001_11110_00010_00000_00001_00000_11111_00000_11111_00001_00000_00010_00000_00001;

		#2
		WriteAddressSelect <= 10'b11100000;  //node 224
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11111_11111_00001_00000_11111_00000_00000_11111_00001_00010_11111_00010_00000_00000_11110_00001_00001_00000_11111_11111_00000_00000_11111_00000_00001_11111_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b11100001;  //node 225
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11110_00000_00001_11111_00000_00010_00000_11111_00000_00001_00000_00000_00000_00001_00001_00000_00000_00000_00001_00000_00000_00001_11110_00000_00000_11110_00001_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b11100010;  //node 226
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11111_11111_00000_11111_00000_11111_00010_00001_00001_00010_11111_00000_00010_00001_00000_00001_11111_00000_00000_11110_00000_11111_00000_00000_00010_11111_00000_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b11100011;  //node 227
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11111_00000_11111_00001_00000_11111_00000_00001_11111_11111_11111_00000_00000_00000_11111_00000_11111_11111_00000_11111_00000_00000_00000_00010_00000_00000_00001_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b11100100;  //node 228
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_00001_11111_11111_11111_11111_00001_00000_11110_11111_11111_00000_11111_00000_00000_00001_11111_00000_00001_00000_00010_00000_11111_00010_00000_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b11100101;  //node 229
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_11111_00000_11111_00000_00000_11111_00001_00001_00000_00001_00000_00001_00000_00000_00000_00010_00000_11111_00000_00000_00000_11110_00000_11111_11111_11110_00000_00000_00001_00010;

		#2
		WriteAddressSelect <= 10'b11100110;  //node 230
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00000_00010_11111_11111_00001_00000_00000_00001_11111_00001_00010_11111_00010_11111_11111_11111_00001_11110_00001_11110_11111_00001_00000_00001_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b11100111;  //node 231
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00010_00000_00000_00001_00000_00001_00000_00000_00001_00001_11111_00001_00010_00000_00010_00001_00000_00010_00001_00000_00001_00000_00000_00000_00000_11111_11110_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b11101000;  //node 232
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00001_00000_00000_00001_00010_11111_00010_00000_00000_00010_11110_00010_11111_00001_00010_00000_00000_11111_11111_00001_11111_11111_11111_11111_00000_11111_11111_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b11101001;  //node 233
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00010_00000_00000_00001_00000_00000_00000_11110_00001_00001_00001_00010_00010_00000_00011_00000_00000_00000_00001_00000_00000_00000_11101_11111_00000_11111_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b11101010;  //node 234
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11110_11111_00000_00010_11111_00001_00010_11111_11111_00010_00001_00000_00001_11111_00001_00010_00000_00000_00001_00000_11111_11110_00000_00000_11101_11111_00001_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b11101011;  //node 235
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_00000_00001_00000_00000_00001_00000_00001_00000_00001_11111_00000_00000_00000_00010_11100_11111_00000_00000_00001_00000_00001_00000_00000_11110_00000_11110_00000_00010_11111;

		#2
		WriteAddressSelect <= 10'b11101100;  //node 236
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00010_00000_00001_00000_00000_00010_00001_11111_00010_00010_11111_11110_11111_11110_00000_11001_00000_00010_00000_00000_00000_11110_00000_00001_11111_00000_11111_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b11101101;  //node 237
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00010_00001_00010_11111_00000_00010_00001_11111_00000_11110_11111_11110_00000_00000_00001_11010_00000_00000_00010_00001_00000_11111_00000_00010_00010_11110_00001_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b11101110;  //node 238
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11110_11111_00001_00000_00000_00001_11111_00001_00001_11110_11111_11110_11111_11111_00000_11111_11110_00000_11111_00000_00001_00000_00000_00010_00000_00001_00000_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b11101111;  //node 239
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11111_00010_11110_00010_00001_00001_11111_00010_11110_00100_11110_11110_00000_11111_00001_00001_11111_00001_00000_00000_00010_00001_00001_00000_11111_11111_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b11110000;  //node 240
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00001_00010_11111_11110_00001_00100_11110_11111_11111_11110_11111_11111_00000_11110_00001_11111_11111_11111_00010_00001_00010_00010_00000_11110_00000_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b11110001;  //node 241
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11101_00001_00000_00000_00000_11111_11111_00000_00010_11110_11111_11111_00000_00001_11111_11111_11111_00001_00001_11111_00001_00000_00010_00101_00010_00000_11110_00000_11110_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b11110010;  //node 242
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_11111_11111_11110_00000_00000_11110_11100_00000_11111_00000_11111_00000_11111_00000_00001_00000_11110_00000_11111_00000_00000_00001_00001_11110_00001_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b11110011;  //node 243
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11111_00000_00000_11111_00001_00000_00001_11111_11101_11111_11110_00010_11111_00001_11110_11111_00000_00001_00000_00000_00000_00001_00000_00001_11111_00000_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b11110100;  //node 244
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_00001_00000_00001_00001_11011_11111_00001_00000_11111_11111_00010_11111_11110_11110_11110_11111_00001_00001_11110_11110_00000_11111_00000_11110_11110_00001_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b11110101;  //node 245
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00010_11111_00000_00001_11111_11111_00010_11111_00001_00000_00010_11111_00001_00000_00000_11111_00001_00000_11110_11111_11111_11111_00000_00001_00010_00001_00001_00001_11110;

		#2
		WriteAddressSelect <= 10'b11110110;  //node 246
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_11111_00001_11111_00001_00000_00001_00001_00010_00001_00001_00001_00001_00001_00010_11111_00001_11111_00000_00001_11111_11111_00000_00001_00001_11111_00000_00001_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b11110111;  //node 247
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_00000_11111_11111_00000_11111_00010_00010_00001_00000_00001_00010_00001_00010_11111_00001_00000_00000_00000_00000_00000_11111_00001_00001_11111_00000_11111_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b11111000;  //node 248
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00010_00000_11111_00001_11110_11111_00001_00001_11111_00000_11111_00000_11111_11110_00000_00001_00000_00000_00000_00010_00000_11110_11111_00001_00001_00000_11110_00000_00010;

		#2
		WriteAddressSelect <= 10'b11111001;  //node 249
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_11111_00001_00001_00010_00010_11111_00000_00010_00000_00001_00000_11111_00010_11111_11111_00010_00000_00000_00001_00001_00001_00001_11111_11111_00000_00001_00000_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b11111010;  //node 250
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_11110_00000_00000_00001_00000_00000_00010_00000_00000_11111_00000_11111_00000_00000_00001_11111_00000_11111_11111_11111_11111_00001_11111_00000_11110_00000_11111_00010_00010;

		#2
		WriteAddressSelect <= 10'b11111011;  //node 251
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00010_11111_11110_00000_00000_00000_00000_11111_11111_00001_00000_11111_00000_00000_00010_00000_00000_00000_00000_00001_11111_00001_00000_00000_00000_11111_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b11111100;  //node 252
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_11111_11111_00001_00000_00000_11111_00000_00000_11111_00000_11110_11111_11111_00001_00000_11110_00001_00000_11111_00001_00000_11111_00000_00000_00000_11111_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b11111101;  //node 253
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_11111_00000_11111_00001_11110_00000_00000_00000_00001_00000_11111_11111_11111_11111_11111_00001_00001_00000_00001_00010_00000_00001_11111_00000_11111_00000_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b11111110;  //node 254
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00000_00001_00000_00010_11111_11110_00001_00000_00000_11110_00001_00000_00001_00000_00001_00001_00000_11111_11111_11111_00001_11111_11111_00000_11111_00000_00000_11111_00001_00010;

		#2
		WriteAddressSelect <= 10'b11111111;  //node 255
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11111_00001_11111_00000_00000_00001_00001_11111_11110_00000_11110_00001_00001_00000_00000_00001_11111_00001_00000_00001_00000_11111_11111_11111_00000_00001_00001_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b100000000;  //node 256
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00001_11110_00000_11110_00010_11110_00001_00001_00001_11110_11111_00000_00001_00010_11111_00000_00001_00000_00000_11111_11111_00000_00000_00000_00001_00001_11110_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b100000001;  //node 257
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_11111_00000_00001_11110_11111_00000_00010_00001_11111_00000_00000_11111_00010_00001_00000_00000_00001_11111_00001_00001_00001_00000_11111_11110_00000_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b100000010;  //node 258
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_00000_11111_00000_00000_11111_11111_00000_11111_00010_11111_00000_00010_00010_00010_00001_11110_00010_00000_00000_00000_00010_00001_00000_00001_11110_11110_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b100000011;  //node 259
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_00001_00001_11110_00001_11110_11110_00001_00000_00001_00001_11111_00011_00000_00010_00001_00010_11110_00001_00001_11111_00000_00010_11110_00000_11111_00001_11111_11110_00001_00001;

		#2
		WriteAddressSelect <= 10'b100000100;  //node 260
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_11110_00001_11111_00001_00000_00011_00001_00000_00010_11111_00010_00010_11111_00011_00001_00001_11110_00000_11111_00001_00000_00000_00000_00000_00001_11110_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b100000101;  //node 261
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11111_00001_11110_00001_11110_00001_11110_00000_00001_11111_00010_00010_11110_00011_00001_00000_00001_11110_11111_00010_00001_11110_11111_11111_00010_11110_00000_00100_00000;

		#2
		WriteAddressSelect <= 10'b100000110;  //node 262
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_11111_00001_00000_11111_00010_00010_11111_00000_00011_11110_00010_00000_00000_00010_11110_00000_00010_11111_11111_11111_11111_11110_11111_11100_00000_11110_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b100000111;  //node 263
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00000_00001_00000_00010_00010_00000_11111_00010_11110_11110_11110_00000_00010_11011_11111_00001_00000_00001_00001_00001_00001_00000_11110_11111_11110_00010_00000_00000;

		#2
		WriteAddressSelect <= 10'b100001000;  //node 264
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11111_00000_00010_00000_11111_00001_00001_00000_00001_00000_00000_11111_00000_00001_00001_10101_00000_00001_00000_00000_00001_11111_11110_00000_00000_00001_00001_00000_11110_00001;

		#2
		WriteAddressSelect <= 10'b100001001;  //node 265
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_11111_00001_00001_00000_00001_00010_00010_00001_11110_00001_00000_00001_00001_00000_11110_11110_00000_00001_00010_00010_11111_00001_11111_00000_00000_11111_00001_11111_11110;

		#2
		WriteAddressSelect <= 10'b100001010;  //node 266
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_11111_00000_00010_11111_00000_00010_00000_11111_00011_11110_00001_11101_11110_11110_00000_00011_11111_00000_00000_00001_00001_11110_00010_00010_00010_00001_00000_11111_11111_00010;

		#2
		WriteAddressSelect <= 10'b100001011;  //node 267
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00001_11101_11101_00001_00010_11110_00100_11110_00001_00001_00000_11111_11111_00001_00000_00000_11111_00001_00000_11110_00000_00001_00001_11111_11111_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b100001100;  //node 268
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11111_11110_00001_00001_11111_00001_00001_11110_00010_11111_11110_00000_11110_00001_11111_00001_11110_00000_11111_00000_00010_00010_00010_00001_00000_00000_11110_00001_00001_00010;

		#2
		WriteAddressSelect <= 10'b100001101;  //node 269
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_00001_00000_11111_11111_00000_00010_11010_11110_11110_11111_00000_11110_00001_00000_00000_00010_00001_11110_11111_00001_00100_00000_00000_11111_11110_11111_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b100001110;  //node 270
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00010_00000_00001_11110_00000_00010_11101_11011_11111_00000_00000_11111_00001_00000_00000_00000_11111_00001_00000_11111_00100_00001_00001_11111_11110_00001_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b100001111;  //node 271
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_00010_11110_00000_00000_11110_11110_11111_11110_11111_00000_00010_11111_11111_00000_00001_00001_11111_11111_11111_11111_00011_11111_00000_11110_00000_00001_00010_00000_11111;

		#2
		WriteAddressSelect <= 10'b100010000;  //node 272
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00001_00001_11111_00001_00000_11110_11111_00001_11111_11111_11110_00000_11111_00000_11111_11110_00001_00001_00010_11111_11111_00000_00000_00001_00000_00001_00001_11110_00000_00000;

		#2
		WriteAddressSelect <= 10'b100010001;  //node 273
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00001_00000_11111_00001_11110_00000_00010_00010_11111_00000_00001_00001_00001_00000_00000_00000_00001_00000_00000_11110_11111_00010_00001_00000_00001_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b100010010;  //node 274
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11111_00001_11111_00001_11110_11111_11111_00010_00000_11110_11111_00000_00010_00001_11111_11111_11111_11110_00001_00000_00000_11110_00000_00010_11111_00001_00000_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b100010011;  //node 275
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00000_11111_00001_00001_11111_00010_00010_11111_11111_00010_11111_00010_00000_00000_11111_00010_11111_00000_00000_11110_00001_00000_00000_00010_00000_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b100010100;  //node 276
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00001_00001_00001_11111_00000_11110_00000_00010_00000_00000_00001_00000_00001_00000_00000_00000_11111_00000_00010_00001_00010_00000_00001_00000_11111_00010_11110_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b100010101;  //node 277
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_11111_00000_00001_00010_00001_00000_00000_11111_00000_00000_11111_00010_00001_00000_00001_11111_00001_00001_00001_00001_11111_11110_00000_00000_00001_00010_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b100010110;  //node 278
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_00001_11111_11111_11110_00000_00000_11110_00000_00001_00000_11111_00010_11111_11111_00000_00000_00000_00000_11111_00001_00010_00000_00010_00001_00000_11111_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b100010111;  //node 279
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_11111_11111_00000_00000_11111_11111_11111_00000_00000_00010_11111_11110_00000_00000_11110_11111_11111_00001_00010_00000_11111_00001_11110_00000_00001_00000_11111_11111_11111;

		#2
		WriteAddressSelect <= 10'b100011000;  //node 280
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00001_00001_11110_00000_11111_11111_11111_00000_11111_11111_11110_00000_00001_11111_00000_00001_00000_00001_11111_00000_00000_11111_11111_00001_00000_00000_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b100011001;  //node 281
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00010_00001_00000_00001_11111_11111_00000_00000_00001_00000_00000_11111_11111_00000_11111_00000_00000_00010_00000_00001_00000_00000_00000_00010_00000_11111_11110_00001_00010;

		#2
		WriteAddressSelect <= 10'b100011010;  //node 282
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_11110_11110_11110_11110_00000_00001_11111_00000_11111_00000_00001_11111_11111_00000_11111_00000_00010_00001_00000_00000_00000_00000_00000_00001_00001_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b100011011;  //node 283
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00000_00000_00000_11111_11111_11111_00001_00010_00001_00001_00000_00000_00000_11111_00000_11111_00000_11111_00001_11111_11111_00000_00000_00010_00001_11111_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b100011100;  //node 284
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_11111_11111_00000_00001_11110_11110_00001_00001_11110_11111_00001_00000_11111_00000_00010_00000_11110_00000_00000_00001_11111_11111_00000_00000_00001_00000_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b100011101;  //node 285
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_11111_00010_00000_00000_00000_00001_00001_11111_00000_11111_00000_00000_00000_00010_00000_11111_00010_00001_00001_00001_00001_00001_00000_00000_00001_00000_11110_00001_00010;

		#2
		WriteAddressSelect <= 10'b100011110;  //node 286
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_11111_11111_00001_00000_00010_00001_00001_00001_11111_00010_11110_00001_00001_00010_00010_00010_11111_11111_11111_11111_11110_11110_11110_11111_00001_00001_11110_00010_00010_00010;

		#2
		WriteAddressSelect <= 10'b100011111;  //node 287
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00000_00000_11111_11111_11111_00001_00000_00010_00001_00001_00010_00001_00001_00010_00010_11111_00000_00001_00000_00000_00001_11111_11111_00000_00000_11110_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b100100000;  //node 288
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11110_11111_00000_11111_00000_00001_00000_11111_00010_11110_00001_00001_00000_00011_00001_00001_11111_00000_11111_00000_11101_11111_00000_11111_00000_00000_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b100100001;  //node 289
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11110_11110_11110_00001_00001_11111_00001_00010_00000_11111_00010_00000_00010_00000_11111_00011_00000_00000_00000_11111_11111_00000_11111_11101_00000_11110_00000_00000_11111_00010_11110;

		#2
		WriteAddressSelect <= 10'b100100010;  //node 290
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_11111_00001_11111_00001_00000_00010_00010_00000_00000_00010_11110_00010_11111_00000_00100_11110_11111_00000_11110_00010_00001_00001_11111_11111_11010_00001_11110_11110_00001_11111;

		#2
		WriteAddressSelect <= 10'b100100011;  //node 291
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00001_11111_00000_00001_00010_00001_00010_00010_11111_00010_00010_11110_11111_00000_00010_11000_00001_00000_00001_00000_00001_00010_00000_11111_00001_11111_11110_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b100100100;  //node 292
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_11111_00000_00001_00001_00001_00001_00001_00000_00000_00000_11111_00001_11111_00001_11011_00010_00000_11110_00010_00001_11110_00001_00010_00010_00001_00000_11111_11101_00000;

		#2
		WriteAddressSelect <= 10'b100100101;  //node 293
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00000_00000_00001_00000_11110_00010_00001_00001_00010_11110_11111_11110_11111_00000_00001_00000_00000_00001_00000_00001_00001_00010_00010_00001_00011_11110_00000_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b100100110;  //node 294
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_11111_00001_11111_11110_00010_00001_11110_00010_00000_11111_00000_11111_00000_11110_00010_00000_00001_00001_00001_00000_11101_00001_11111_00010_00000_00000_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b100100111;  //node 295
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_00001_11111_11101_00010_00001_11111_00011_11111_00000_00000_11111_00000_11111_00010_00001_00001_11110_00000_00000_11110_00001_11110_00010_00001_11110_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b100101000;  //node 296
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00010_00000_00000_11110_00000_00001_11111_00011_00000_00001_11111_11101_00000_00000_00000_11111_11111_11110_00001_00001_00010_00010_11110_00000_11110_11110_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b100101001;  //node 297
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00000_00001_00000_00000_11110_00010_00010_11011_00010_11111_00000_00000_11101_00010_11110_00000_11111_00001_11111_00000_00000_00011_00000_00000_00001_00000_00000_00010_00001_11111;

		#2
		WriteAddressSelect <= 10'b100101010;  //node 298
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00010_00000_00001_11110_00001_00000_11110_11110_11110_11110_00001_11110_00010_00001_11111_00001_00001_00000_00001_00000_00010_11111_00010_11111_11101_00001_00001_00010_00001;

		#2
		WriteAddressSelect <= 10'b100101011;  //node 299
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11110_00010_11101_00000_11111_11110_00010_11111_11100_11110_11110_00000_00001_00000_11111_00000_00001_11111_00000_11111_11110_00001_11110_00001_11110_11111_00010_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b100101100;  //node 300
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00010_00000_11111_00000_11110_00001_00010_11110_11111_00000_00010_00001_11111_11111_11111_00001_00001_11111_00000_00000_00000_00001_00010_11110_11111_00010_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b100101101;  //node 301
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_11110_00000_11111_11110_11111_11111_00001_00001_00000_00001_00001_11111_00001_00001_00010_00010_00000_11110_00001_11111_00000_11111_00000_00001_00000_11111_00000_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b100101110;  //node 302
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00000_00010_11111_11110_11111_00000_00010_00010_00000_00000_00000_00001_00001_00010_11110_11110_00000_11110_00000_00001_00000_11110_00010_00000_00000_00000_00001_00001_11110_00001;

		#2
		WriteAddressSelect <= 10'b100101111;  //node 303
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_00010_00001_11111_11111_11111_11110_00010_11111_00000_00000_00010_11111_00010_00000_00000_00001_00010_11110_00000_00000_11111_00001_00010_00000_11111_00001_11110_00010_11111;

		#2
		WriteAddressSelect <= 10'b100110000;  //node 304
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_00010_00001_00000_00000_00001_00000_00000_00010_00000_11111_11111_00000_00001_00000_11110_00001_00001_00001_00000_00000_00001_11110_00000_11111_11111_11111_00000_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b100110001;  //node 305
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_11111_00000_11110_00001_00010_00000_00001_11110_11111_00001_00000_11111_00010_00000_00010_11111_00000_00001_11110_00000_00010_00000_11111_11111_00000_00001_00000_00000_00001_00010;

		#2
		WriteAddressSelect <= 10'b100110010;  //node 306
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_00001_00000_00010_00001_00000_11111_11111_11111_00000_00001_11111_00001_11111_00000_11111_11111_00000_00000_11111_00001_00001_11111_00000_00001_11111_11111_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b100110011;  //node 307
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00010_00001_11111_00001_00001_00010_11111_11111_00000_11111_11110_00000_00000_00000_11111_00000_00000_11110_00000_11111_11111_00000_11110_00000_00000_00000_11110_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b100110100;  //node 308
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11111_00000_00000_11111_00000_00001_00001_00000_00001_00000_11111_00010_00000_11110_00010_00010_00000_11111_00001_00010_00001_00010_00000_00000_11111_00001_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b100110101;  //node 309
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11110_11111_00001_00001_11111_00000_00010_00010_00001_00000_00001_00000_11111_11110_00000_00000_00000_00000_11111_11110_11111_00001_11111_00000_00000_00001_00000_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b100110110;  //node 310
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_00001_11111_00000_00000_00000_11111_00000_00001_11111_00000_00001_00000_00000_00000_11111_00000_00000_00000_00000_00000_11111_00001_00000_00000_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b100110111;  //node 311
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00000_00000_11111_11111_00000_11110_11110_00000_11111_00000_00001_00000_00001_00000_11110_00001_11111_11110_00001_11111_11111_11111_11111_00010_00000_00001_00000_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b100111000;  //node 312
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11110_11111_11110_00010_00001_00001_00010_11111_11111_11110_00010_00000_11111_00001_00000_11110_00001_00000_00000_11111_00000_00010_00000_11111_00010_11110_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b100111001;  //node 313
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_11111_00001_11111_11110_00000_00001_00000_11111_11110_11111_00001_00000_00001_00001_11110_00000_00010_11111_11110_11110_00010_11111_00000_00000_11110_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b100111010;  //node 314
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_00000_00000_00000_11111_00000_11111_00010_00000_11111_00000_00000_00000_00010_00001_00000_11111_00001_11111_00010_11110_11111_00000_11110_00001_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b100111011;  //node 315
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_00001_00001_11110_11110_11111_00001_00000_11111_00000_00000_00010_11111_00000_11110_00010_11111_00001_11111_11111_00000_00000_11110_11111_11111_00010_00000_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b100111100;  //node 316
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11100_00000_00010_11111_11111_00000_00010_00000_00001_00010_00001_00001_11111_11110_11110_00011_00001_00010_00010_00000_00000_11110_00010_11111_11110_11111_11110_11110_00001_00001;

		#2
		WriteAddressSelect <= 10'b100111101;  //node 317
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00010_00001_00001_00000_11111_00001_00000_11110_00010_00000_00010_00010_11111_00001_00000_11110_00010_11110_00010_00001_00010_11111_11111_11110_00010_11110_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b100111110;  //node 318
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00010_00000_00010_00010_11111_00000_00010_00000_11111_00010_00000_00100_11110_11111_00001_11101_00001_00010_11110_00001_00000_11111_11111_11111_11101_00100_00000_11111_00010_00001;

		#2
		WriteAddressSelect <= 10'b100111111;  //node 319
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00010_11110_00001_00001_00000_00000_00010_00001_11110_00011_00000_00001_00000_11111_00010_11010_00001_00001_11111_00010_00000_11110_00001_00000_00000_11111_11110_11110_11111_11110;

		#2
		WriteAddressSelect <= 10'b101000000;  //node 320
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00010_00010_00010_00001_00010_00010_00001_11111_11110_11110_11111_11110_00010_00000_00000_11110_00010_00001_00010_00010_00001_11110_00000_00001_00010_00001_00000_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b101000001;  //node 321
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_11111_00010_11111_11111_00010_11111_00001_11111_11110_11111_11110_00001_00000_00001_00000_00000_00001_00000_00010_00001_00000_00010_00000_00100_00000_11111_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b101000010;  //node 322
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_00000_00000_11111_00000_11110_00010_00000_00000_00000_11110_11111_11101_00000_00001_11110_00001_00001_00001_00000_00000_00010_11110_00010_11111_00010_11110_11110_00000_00010_11111;

		#2
		WriteAddressSelect <= 10'b101000011;  //node 323
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11111_00000_00010_00001_11110_00010_00000_00000_00100_11110_11110_11111_00010_00000_11111_00010_11111_00000_00010_00000_00001_11110_00010_00000_00010_11111_11110_00010_11110_11111;

		#2
		WriteAddressSelect <= 10'b101000100;  //node 324
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_00011_00001_00001_11110_00010_00001_00000_00101_11110_11110_00001_11110_00000_11110_00001_00000_00001_11111_00001_00001_00010_00001_00000_00000_11111_11110_00010_00000_11111;

		#2
		WriteAddressSelect <= 10'b101000101;  //node 325
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00001_11110_00010_11111_00000_00000_11011_00010_11111_00000_00010_11011_00001_00000_00010_11111_00001_00010_00010_00000_00010_00010_11111_00010_11110_11110_00010_00001_11111;

		#2
		WriteAddressSelect <= 10'b101000110;  //node 326
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00010_11110_11111_11110_00000_00010_11010_00001_11110_11111_00001_11110_11110_11111_00000_00001_00000_00001_00000_11111_00011_00001_00001_00001_11101_00000_00010_00001_00001;

		#2
		WriteAddressSelect <= 10'b101000111;  //node 327
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_00000_11110_11110_11110_11110_11111_11111_11010_11110_00001_11111_00000_11111_00000_00000_00001_11111_00010_00000_11111_00011_00010_00010_11111_11110_00000_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b101001000;  //node 328
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_00010_11110_11110_11111_11111_00000_00001_11111_11111_00001_00010_00001_11110_00010_00000_00001_11100_00000_11110_00000_11110_00001_00000_11111_00000_00010_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b101001001;  //node 329
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00001_00000_00001_00001_11111_00001_00100_11110_00000_11111_00001_00001_00010_00000_00000_00000_00000_00000_11111_11111_11111_00001_00001_00000_11111_00000_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b101001010;  //node 330
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00001_00000_00001_00001_00001_00000_00010_00011_00000_00000_00001_00001_00000_00010_11111_11111_00010_00010_11110_00000_00001_11111_00010_00010_11111_00000_00010_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b101001011;  //node 331
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_11111_00000_00001_11111_11111_00001_00000_00010_00010_00001_11111_00010_00010_00010_11111_00001_00000_00000_11111_11110_00001_00001_00010_00001_00010_11110_11111_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b101001100;  //node 332
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_00000_00001_00001_11110_00000_11111_00000_00001_00001_00000_11111_00000_00001_00000_11110_00001_11111_00010_00001_11111_00001_11111_00000_00000_00000_11111_11111_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b101001101;  //node 333
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_00000_11111_00010_11111_00000_00001_00001_00010_11111_00010_00000_11111_11110_00001_00000_00000_11111_00001_00001_00000_11111_00010_00000_00001_11111_11110_00001_00010;

		#2
		WriteAddressSelect <= 10'b101001110;  //node 334
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_11111_00010_00000_00000_00000_00000_00000_00001_11111_00000_00001_11111_00000_11111_00001_00001_11111_11111_00001_00001_00000_00000_00001_00000_00001_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b101001111;  //node 335
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00001_11111_00000_11111_00000_00000_11111_00010_00001_11111_00000_00010_00000_11111_11111_00000_00000_00000_00000_00000_00000_11111_00000_11111_00000_00000_11110_00000_00000;

		#2
		WriteAddressSelect <= 10'b101010000;  //node 336
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_11111_11110_00001_00000_00000_00010_00000_00000_00001_00000_00000_00000_11110_00001_00001_11110_00001_00000_00000_00000_00000_00000_00000_00000_00000_00000_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b101010001;  //node 337
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_00001_11111_00010_11111_00000_11111_00000_00000_00001_00000_00000_00010_00000_00000_00000_00000_00000_00001_00001_00000_00000_00010_11111_00010_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b101010010;  //node 338
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00000_11111_00000_00001_00000_00010_11110_11111_00010_00001_00000_11111_00000_11110_11111_00001_00000_00000_00001_00010_00001_11110_00001_11111_00001_11111_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b101010011;  //node 339
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_11111_11111_00000_11111_11111_00001_11110_00010_11110_00000_00010_00000_00000_00000_00001_00000_11111_11111_00000_00000_00000_00010_00000_00001_11110_00000_11111_00010;

		#2
		WriteAddressSelect <= 10'b101010100;  //node 340
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00001_00000_00001_11111_00001_11111_00000_00001_00001_00001_11110_00001_00010_00001_00000_00001_11111_00000_00000_00000_11110_00000_00001_00000_00000_00000_00000_11111_11111_11111;

		#2
		WriteAddressSelect <= 10'b101010101;  //node 341
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11110_00000_00000_00001_00001_00001_11111_00000_00000_11110_11111_11111_00010_00010_11111_00000_11110_11111_00001_11110_00000_00001_00000_11111_00001_00000_11110_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b101010110;  //node 342
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00001_00000_00010_00001_11111_00000_00001_00010_00001_00001_11111_00001_00001_00010_11111_00010_11111_00011_00001_11111_11111_00010_00001_11111_00011_00000_11111_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b101010111;  //node 343
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11110_11110_00001_11110_11111_11111_00010_00000_11111_00010_00000_00001_00001_00000_11010_11111_00000_00001_00001_00000_00000_00010_00001_00000_00000_00001_11111_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b101011000;  //node 344
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00010_00010_11111_00000_00000_00010_00000_00001_00001_00001_00101_11110_00001_11100_11111_11110_00010_11111_00000_00010_00000_11110_11111_11110_00010_11110_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b101011001;  //node 345
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_11111_00010_00001_00001_11110_00000_00000_00000_11110_00010_00010_00011_11111_11110_11101_00001_11111_00001_00000_00000_00100_00010_00000_11110_11101_00001_11111_11110_00001_11111;

		#2
		WriteAddressSelect <= 10'b101011010;  //node 346
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00010_00001_00001_11111_00001_00000_00000_00001_00001_00000_00011_00000_11111_11110_11010_11110_00000_11111_00010_00001_00000_11110_00000_11110_00010_00000_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b101011011;  //node 347
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00100_00010_00010_00001_00010_00000_11111_00001_00000_00010_00000_00001_00011_11111_00000_11010_00011_00001_00001_00010_00001_00000_00001_11110_00011_00001_11111_00000_11110_00001;

		#2
		WriteAddressSelect <= 10'b101011100;  //node 348
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00010_00000_00010_00000_00010_00000_11110_00000_11111_11110_00000_11110_00001_00000_11111_11111_00001_00010_00000_00001_11110_11111_00010_00001_00101_00001_11111_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b101011101;  //node 349
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00000_00000_00000_11110_00001_00010_11110_11110_11111_11110_00001_11111_00010_11111_11111_00000_00010_00011_00000_00010_11101_11111_00010_00000_00011_00000_00010_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b101011110;  //node 350
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_11111_00000_00000_00000_00000_00001_11110_00001_00000_11110_11110_11110_00010_11111_11111_00010_00001_00000_11101_00000_11111_11110_00001_11111_00010_11111_11111_00010_00000_00000;

		#2
		WriteAddressSelect <= 10'b101011111;  //node 351
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_00000_00000_00000_00011_11111_00000_00101_11110_00000_11111_11110_00010_11111_00010_00000_00001_11111_11111_00000_11110_00010_11111_00001_11111_00010_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b101100000;  //node 352
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00010_00000_00001_11111_00010_11111_00001_00100_00000_11110_00000_11111_00010_00000_11111_00000_00010_11111_00001_11111_11110_00010_00001_00010_00000_00000_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b101100001;  //node 353
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11110_00010_11110_00010_11110_00001_11111_11101_00011_11101_00000_00001_11101_00000_00000_00000_00000_00000_11111_00010_00010_00010_00001_00001_11111_11110_11111_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b101100010;  //node 354
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_00010_11101_11111_11111_00001_00000_11010_00000_11111_00001_00010_11100_00001_11110_00000_00000_00010_00000_11111_00000_00010_00001_11110_00001_11100_00000_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b101100011;  //node 355
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_00001_11110_00001_11111_11101_00010_11110_11110_11101_00010_00001_11111_00000_00001_00000_00000_00001_00001_00000_00000_00010_11110_00001_00000_11011_00000_00010_00000_00001;

		#2
		WriteAddressSelect <= 10'b101100100;  //node 356
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_11111_11111_11111_00001_11110_11110_00001_00000_11110_11111_00010_00000_11111_00001_00001_00000_11111_11111_11111_00000_00000_00000_11111_00001_11111_11111_00010_00010_11111_00001;

		#2
		WriteAddressSelect <= 10'b101100101;  //node 357
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00001_00000_00001_00000_11111_00001_00100_11110_00000_00000_00000_11110_00010_00001_11111_00001_11111_00001_11111_11111_11111_00001_11110_00000_00000_00010_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b101100110;  //node 358
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00000_00010_11111_00001_11110_00000_00010_00010_00001_11111_11111_00001_00011_11111_00000_11111_00001_00001_11111_11111_00001_00001_00001_00000_00001_00001_00010_11110_11111;

		#2
		WriteAddressSelect <= 10'b101100111;  //node 359
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00000_11111_11111_11111_00000_00001_00010_00001_00000_00000_00010_00001_11110_00010_00001_00001_11110_00010_11110_00000_11111_00000_00010_00001_00001_00010_00000_00001_00010_00001;

		#2
		WriteAddressSelect <= 10'b101101000;  //node 360
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00000_00000_00000_11111_11110_00001_00010_00001_11111_00000_00010_00010_00001_00000_11111_00001_00010_11111_11111_00001_11111_00000_00010_00000_00000_00000_00010_00000_00001;

		#2
		WriteAddressSelect <= 10'b101101001;  //node 361
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00000_00000_00000_00010_11110_00001_00001_00000_00001_11111_00000_00000_00001_11111_00001_00001_00001_11111_00001_11111_00000_11111_00000_00000_00000_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b101101010;  //node 362
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11110_11111_11111_11111_11111_00010_00000_11110_00000_00000_00010_11110_00001_00000_00000_11111_11111_00010_11110_00001_00000_00000_00000_00010_11110_00000_11110_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b101101011;  //node 363
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00001_00000_11110_11111_00000_11111_00000_00001_00000_00001_00000_11111_00000_00001_00001_00000_11111_00000_00000_00000_00001_11111_00000_11111_11110_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b101101100;  //node 364
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_11111_00000_00000_11111_00001_11111_11111_00001_11111_00001_00001_00000_00010_00001_00000_11111_00001_11111_00000_11110_00000_00000_00000_00001_00000_00001_00000_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b101101101;  //node 365
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00001_00001_00000_00000_00001_11111_11110_00001_00000_11111_11111_00001_00001_11111_00000_00000_00001_00000_00000_11111_11110_11111_11111_00001_00001_11111_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b101101110;  //node 366
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00001_00000_00000_11110_00001_00000_00000_00000_11111_00001_00000_00001_00000_00001_00000_00001_00001_11110_11111_00000_00000_11110_11111_00010_11111_00001_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b101101111;  //node 367
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_00001_00000_00000_00001_11111_11110_00000_00001_00001_00000_11111_11111_00001_00001_00000_00001_00001_11111_00001_00001_00001_11111_11111_00001_00001_00000_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b101110000;  //node 368
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00000_11111_00000_00001_11110_11111_00000_11111_11111_00001_00000_00001_00001_11111_00001_11111_00000_00000_11111_00000_11111_00000_00000_00000_00010_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b101110001;  //node 369
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00000_00000_11110_00000_11111_00001_00001_11111_00000_00000_00000_00001_00010_11100_00010_11111_11111_00001_11110_00000_00000_00001_00001_00000_00010_11110_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b101110010;  //node 370
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_11111_11111_11110_00010_11111_00000_11111_11111_11111_00000_11111_00010_00000_00001_11100_00001_00000_11111_00001_11110_00001_11111_00000_00000_00000_00010_00001_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b101110011;  //node 371
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11101_00000_11111_00000_11110_11111_11111_00010_11111_11111_11111_00001_00001_00001_11010_00010_00010_11110_00000_11111_00000_11111_00001_00000_11111_00010_11110_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b101110100;  //node 372
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11111_00001_00000_00000_00000_00000_00000_00000_00000_11111_00001_00010_00000_00001_11010_00010_00001_00000_00000_00000_00010_00000_00000_11101_00000_00000_00000_11110_00010_11110;

		#2
		WriteAddressSelect <= 10'b101110101;  //node 373
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00010_00001_00000_00000_11111_00001_00001_00010_00000_11111_00000_00011_00000_00000_11011_11111_11111_11111_11100_00001_00010_00001_00001_00000_11110_00011_11111_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b101110110;  //node 374
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00010_00010_11110_00000_00010_00001_00010_11111_11111_00011_00001_00100_11110_11111_11100_11011_11111_11111_11111_00010_11111_00001_11111_11110_00010_00010_00010_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b101110111;  //node 375
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00010_00000_11110_11110_00000_11110_11111_00000_11110_00010_00010_00001_00010_00000_11111_11100_11110_00001_00010_00000_11110_11110_00000_11111_00101_00000_00010_00010_00000_00001;

		#2
		WriteAddressSelect <= 10'b101111000;  //node 376
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00011_00000_00000_00010_00000_11110_00010_00010_11101_00001_00000_11101_00001_11111_00001_00000_11111_00000_00010_00000_00000_00010_00001_11110_00001_00000_00011_11111_00000_00010_00010_11111;

		#2
		WriteAddressSelect <= 10'b101111001;  //node 377
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00010_00010_11111_11111_00010_00010_11110_11111_00000_11110_11111_11111_00010_11111_11110_00001_00010_00000_00000_00001_11111_00000_00001_11110_00010_11110_11110_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b101111010;  //node 378
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_11110_00010_11110_00001_00001_00010_11110_11111_00000_00000_00000_11110_00011_00001_00000_00010_00010_00000_00000_00000_00000_11110_00000_11111_11110_11111_00000_00001_00000_11110;

		#2
		WriteAddressSelect <= 10'b101111011;  //node 379
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00011_11111_00010_00010_00000_11110_00000_00010_00000_00000_11111_00010_11111_00001_00010_00000_00000_00001_11101_00000_00000_00010_11101_11111_00001_00001_00010_00010_00001;

		#2
		WriteAddressSelect <= 10'b101111100;  //node 380
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00011_11110_00000_00010_11101_00010_00010_11111_11101_00000_00010_11110_00010_00001_00000_00010_00000_00010_00010_00010_00001_11111_00001_00001_00001_11110_00000_11110_11111_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b101111101;  //node 381
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_11111_00001_11110_00010_00010_00001_11111_11110_00010_11111_00010_00001_11011_11111_00000_00001_00010_00001_00000_00010_00000_00010_00010_11111_00001_11110_11101_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b101111110;  //node 382
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11111_11111_11110_00010_00001_00000_00000_11011_00001_00000_00010_11111_11110_11111_00001_00010_00010_00001_00001_11110_00001_00010_00011_11111_00000_11110_00010_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b101111111;  //node 383
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00010_11111_00000_00000_00001_11110_11111_00000_00000_11110_00011_00010_00000_00000_00001_00000_00001_11111_00001_00000_11110_11111_00000_11111_00001_11111_00001_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b110000000;  //node 384
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_11101_00000_00000_11111_11110_00010_00001_00001_00001_11111_00010_00001_00001_00010_00001_00000_11111_00000_00000_00001_00010_00010_11111_00000_00001_00010_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b110000001;  //node 385
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00001_11110_00010_00010_00000_00001_00010_00000_00000_11111_00001_00000_00001_00001_00000_00001_00001_11111_00000_11111_00000_00000_00000_00001_00010_00010_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b110000010;  //node 386
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00000_00000_00001_00000_11111_00001_00010_11111_00000_11111_00001_00000_00010_00001_00000_00000_11111_00000_00000_11110_00001_00001_00000_11111_11111_00001_00001_11111_00010;

		#2
		WriteAddressSelect <= 10'b110000011;  //node 387
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_00000_11111_00000_00010_00001_00000_11111_00010_11111_00000_00000_00001_00010_00011_00001_00001_00000_00010_11111_00000_11111_11111_00001_00001_00001_00000_11111_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b110000100;  //node 388
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00000_00010_11111_00010_00000_00001_00000_00001_00001_00000_00010_00000_00001_00000_00000_00001_00010_00000_00000_00001_00001_00000_00000_00000_11111_11110_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b110000101;  //node 389
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_11111_00000_00000_00010_00000_00000_00000_00001_00010_00000_00000_00001_00000_00000_11111_00000_00010_00010_11111_00000_11111_11110_00001_00001_00000_11110_11110_00010_11111;

		#2
		WriteAddressSelect <= 10'b110000110;  //node 390
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_11111_00010_11111_11111_00001_00001_11111_00000_11110_00000_00001_11110_00000_00010_11111_00000_00000_00001_11111_00000_11110_00001_00000_00000_00001_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b110000111;  //node 391
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00010_00001_00000_00010_11110_00001_00000_11110_00010_00000_11111_00001_00000_11111_00000_11111_00000_00010_00000_00001_00000_00001_00001_00000_00000_00000_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b110001000;  //node 392
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_11110_00001_00000_11111_00000_11110_00000_00001_00001_00000_00001_00010_11111_11111_11111_00000_00000_00010_00001_00010_00000_11111_00000_11111_00001_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b110001001;  //node 393
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_00000_00001_00000_11110_11110_11111_00000_11111_00001_00000_00000_11111_11110_00000_11111_00001_11110_00000_11111_11111_00010_11110_11111_00000_00000_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b110001010;  //node 394
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00010_00000_11110_00000_00001_00010_00001_11111_00001_11111_00000_00001_11111_00000_00000_00000_00000_00000_00001_11111_00000_00010_00000_11111_00000_00000_11111_00001_11110_00001;

		#2
		WriteAddressSelect <= 10'b110001011;  //node 395
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11111_11111_00000_11110_00000_00000_00000_00000_00010_11111_00000_00001_00000_00001_11110_11111_00001_11110_11111_11111_00001_00001_11111_00001_00001_00010_11111_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b110001100;  //node 396
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_00000_11111_11111_00001_11110_11111_11111_00001_00000_11110_11101_00000_00001_00000_00000_00001_11111_11111_11111_11111_00001_11111_00000_11110_00010_11111_00000_00001_11110;

		#2
		WriteAddressSelect <= 10'b110001101;  //node 397
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_11111_00010_00001_00000_00010_00001_00001_11110_00001_11111_00000_00010_11110_00000_11111_00001_00000_00000_11111_00001_00001_00001_11111_00001_11111_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b110001110;  //node 398
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11111_11111_11111_11111_00001_00001_00001_11111_11111_00001_00010_00001_00001_11011_00001_00001_11110_00010_00001_00001_00000_00010_00000_00010_00010_11110_11110_00011_00001;

		#2
		WriteAddressSelect <= 10'b110001111;  //node 399
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11011_00010_11101_00000_00010_11111_11111_00001_11111_00010_00000_11111_11111_00001_11110_00010_00000_11111_00010_00010_00000_00010_00000_11110_00001_00010_00000_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b110010000;  //node 400
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00001_00010_11110_00010_11111_00000_11111_00010_00000_00000_00010_00010_00001_00010_11110_00011_00000_11110_11111_00000_00000_00000_11111_11110_00001_00001_00001_00001_00010_11111;

		#2
		WriteAddressSelect <= 10'b110010001;  //node 401
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_11110_11111_00001_11110_00000_00000_00000_00001_00001_00011_11110_11110_11110_11110_11110_11110_11100_00010_11111_00000_11110_11010_00001_00000_00000_11111_00010_11111;

		#2
		WriteAddressSelect <= 10'b110010010;  //node 402
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00001_11110_11110_00010_11110_00010_00001_11111_00001_00010_00011_11110_11110_11110_11101_11011_11110_11110_00001_11111_11110_11111_11110_00001_00000_00001_00001_00011_00001;

		#2
		WriteAddressSelect <= 10'b110010011;  //node 403
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00010_00010_11101_00000_00011_11110_00001_11111_11101_00010_00010_11110_00001_00000_11110_11111_11110_00001_00010_11111_11101_11101_00001_11110_00010_11110_00001_00010_00000_11111;

		#2
		WriteAddressSelect <= 10'b110010100;  //node 404
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00001_00001_11110_11111_00011_00001_00001_11110_11110_11111_00010_11110_00010_11110_11111_00000_11110_11111_00010_00000_11111_00000_11110_11110_00001_11111_00010_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b110010101;  //node 405
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00000_00001_11101_00010_00010_00001_00000_11111_00000_00001_00010_11111_00010_00010_11111_00001_11111_11110_11111_11111_00001_11101_11110_11110_11110_11111_00001_00001_11110_11110;

		#2
		WriteAddressSelect <= 10'b110010110;  //node 406
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00010_11111_00010_00100_00010_00000_00010_00010_00000_00010_11111_00010_00010_00010_00010_00001_00010_00000_00000_00001_00000_00001_11110_00000_11111_00000_00001_11110_00001;

		#2
		WriteAddressSelect <= 10'b110010111;  //node 407
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00000_00010_11110_00001_00011_00000_11110_00000_00010_00000_00010_11110_00001_00001_11111_00000_00001_11111_11111_00001_00010_11110_00010_11111_11111_00001_11111_00010_11111_11111;

		#2
		WriteAddressSelect <= 10'b110011000;  //node 408
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00001_11111_11110_00001_00010_00000_00001_11111_00001_00000_00010_11111_11110_11111_00001_00010_00001_11110_00000_11111_11111_00000_00010_11111_11111_00001_00000_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b110011001;  //node 409
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00000_11110_00000_00001_00001_00010_00000_11101_00000_00001_00010_00010_11110_11111_11111_00000_00001_11111_00000_11111_00001_00001_00010_00000_00010_00001_00000_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b110011010;  //node 410
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11110_11110_00000_00001_00000_00000_00000_11101_11110_00001_00010_11111_11111_11110_11111_00000_00000_00000_00000_00000_00000_00001_00010_11111_11111_00000_00010_00000_11111_00010;

		#2
		WriteAddressSelect <= 10'b110011011;  //node 411
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11111_11101_00001_11111_11111_11110_00000_11111_11111_00001_00000_00001_11111_00000_00001_00010_00000_11111_11111_11111_00000_00001_00010_11111_00001_00010_00001_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b110011100;  //node 412
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_11111_00000_00001_00000_00010_11110_11111_00000_00001_11111_00001_00000_11111_00000_00001_00000_11111_11111_00001_11111_00000_00000_11111_00001_00000_00000_00010_11111_11111_00010;

		#2
		WriteAddressSelect <= 10'b110011101;  //node 413
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_00000_00001_00001_11101_00001_00010_00000_00000_00000_11111_00001_00110_00010_11111_00001_00000_11111_11111_00000_00000_00000_11111_00000_00001_00001_00001_11111_11110;

		#2
		WriteAddressSelect <= 10'b110011110;  //node 414
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00001_00000_00000_00010_11111_00010_00010_00000_11111_00001_00000_11111_00010_00001_00010_11111_00000_00000_11110_00000_00001_11111_11110_11110_00000_00001_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b110011111;  //node 415
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_11110_00010_00000_00000_11111_00010_00001_00000_11111_11111_00000_11111_00010_00000_11110_00000_00001_11111_00000_00010_00001_11111_00000_00000_00000_00000_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b110100000;  //node 416
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_11110_11111_11111_11111_11111_00001_00001_00001_11111_11110_00010_00000_00000_00001_00000_00000_00001_00000_11111_11111_11111_11110_00000_00010_11110_11110_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b110100001;  //node 417
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00000_00010_00000_11111_11111_00001_00000_00000_00001_11111_00000_00001_00000_00000_11111_11111_00000_00000_00000_00000_11111_00000_11111_00000_00000_11110_11110_00010_00000;

		#2
		WriteAddressSelect <= 10'b110100010;  //node 418
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00010_11111_00000_11111_11111_00001_11111_00000_00010_00000_00000_00001_11111_11111_00000_00001_00000_00000_00001_00001_00000_11111_00010_00000_00010_11110_00000_00010_00010;

		#2
		WriteAddressSelect <= 10'b110100011;  //node 419
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11110_00001_00001_00001_11111_11111_11111_11110_00000_00001_11111_11111_11111_11111_00001_00000_00010_00000_00000_00000_00000_11110_00000_00000_00000_00001_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b110100100;  //node 420
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_00000_00000_11111_11111_00000_11111_00000_00001_00001_11110_00000_00000_11110_11110_00000_00000_00000_00000_11110_00000_11111_00001_11110_00001_00000_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b110100101;  //node 421
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00000_00000_11111_00000_11110_00001_00000_11111_00010_11111_00000_00000_00000_11111_11111_11111_00000_00000_11111_11111_11111_00001_11111_00000_00000_00000_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b110100110;  //node 422
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_00001_00001_11111_11111_11111_00001_00000_00000_00000_00000_00000_00001_00001_00000_00000_11110_11111_00000_11111_00000_11111_00001_11111_00000_00001_00000_00001_11111_11110;

		#2
		WriteAddressSelect <= 10'b110100111;  //node 423
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11111_11111_00001_11111_00000_11111_11111_00000_00001_00000_00000_11111_00001_00010_11110_00001_11111_00001_11111_00000_11111_00001_11111_00010_00000_00001_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b110101000;  //node 424
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_11111_00000_00001_00000_00000_00010_11110_11111_00000_00010_00010_00010_00001_11110_00001_00001_00000_11110_00000_00000_00000_00001_00000_00001_11110_11110_11110_11110;

		#2
		WriteAddressSelect <= 10'b110101001;  //node 425
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_00001_11110_11111_00010_11111_00001_00000_11111_11110_11111_00000_00001_00001_11110_00000_00001_11110_00001_11110_11110_11111_00000_00001_00010_00010_11111_11110_11111_00001;

		#2
		WriteAddressSelect <= 10'b110101010;  //node 426
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_00001_11110_00000_00010_11111_00000_00001_00000_00001_00001_11111_11110_00010_11111_00010_00000_11110_00010_11110_11111_00000_00010_11110_00000_00000_00000_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b110101011;  //node 427
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_11111_11111_00000_00001_11111_00000_00000_00000_11111_00001_00000_00010_00010_00010_11111_00010_11101_00000_00001_00001_00001_00000_11111_00001_00001_00000_00000_00010_00010;

		#2
		WriteAddressSelect <= 10'b110101100;  //node 428
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_11111_00010_00000_00001_00000_00001_00000_00000_00001_00001_00000_00001_11111_00010_00010_00001_00010_11110_11101_00001_00001_00000_00001_11110_00010_00001_11111_11110_00010_00001;

		#2
		WriteAddressSelect <= 10'b110101101;  //node 429
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_00001_11110_00001_00000_11111_11110_11111_00000_00010_00000_00001_00010_11111_00001_00010_11111_11110_11100_00001_00000_00000_11111_11010_00000_00000_00010_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b110101110;  //node 430
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00001_11110_11110_00001_00001_00000_11110_00001_00010_00011_00001_11111_00001_00001_11110_11011_11111_11110_00010_11101_00000_11110_11010_00010_11111_00010_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b110101111;  //node 431
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_00000_11110_00001_00001_11101_11111_11110_11110_00001_00010_11110_00001_11100_00010_00000_11110_00000_00011_00010_00001_11111_00000_11110_00001_11101_00010_11110_00000_11110;

		#2
		WriteAddressSelect <= 10'b110110000;  //node 432
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_00010_11111_00000_00010_00011_00001_00010_11110_11110_00001_00010_00000_00011_00000_00001_00010_00000_00000_00010_00010_00001_00000_11111_11110_00000_00000_00010_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b110110001;  //node 433
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11110_11111_00010_00010_00001_00001_11110_11111_00010_00010_11110_00010_00001_00000_00000_00010_00000_11111_00000_00001_11111_11111_11110_11111_00000_11111_00010_00000_11111;

		#2
		WriteAddressSelect <= 10'b110110010;  //node 434
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_11110_11111_11110_00001_00010_00001_00001_00000_00001_00000_00010_00000_00000_00001_11111_00001_11111_00000_00000_00001_00001_11111_00010_00000_00000_11110_00001_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b110110011;  //node 435
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00000_11100_11110_00010_00010_00001_11110_11101_00010_00001_00010_11101_11110_11111_00000_00001_00001_00000_00010_00000_00000_11111_00010_00000_11111_00001_11111_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b110110100;  //node 436
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_11111_00010_00010_00001_00000_11110_11110_00001_00000_00010_11111_11111_11110_00001_00001_00010_11111_00001_00000_00000_00000_00010_11111_11111_00010_11111_00010_11111_00001;

		#2
		WriteAddressSelect <= 10'b110110101;  //node 437
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_11100_00001_11110_11111_00100_11111_11110_00000_00010_00000_00000_11111_11111_00000_00000_00001_11111_00001_00000_11110_11111_00001_00000_00000_11111_00001_00001_11111_00010;

		#2
		WriteAddressSelect <= 10'b110110110;  //node 438
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_11110_00001_00001_11111_00000_11111_11110_11111_00001_11110_00000_11111_11111_11111_00000_11111_11111_11111_11111_11111_00000_00000_11110_00001_00010_00010_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b110110111;  //node 439
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00011_00000_11110_00010_11110_11111_00000_00000_00000_00000_00001_11110_00000_00000_11101_11111_11111_00000_00000_00000_11111_11110_00001_00001_00001_00000_00010_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b110111000;  //node 440
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11110_11111_11111_00000_00010_11110_00000_00010_00010_00000_00000_00010_00000_00000_00001_00000_11111_00010_00001_00000_00000_00000_00010_00000_00000_00010_11111_00010_11110_00010;

		#2
		WriteAddressSelect <= 10'b110111001;  //node 441
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_11111_11111_00001_11111_11110_00001_00010_00001_00000_11111_00001_00010_00010_00010_11111_00000_00000_00000_11110_11110_00000_00000_00000_11111_00010_00001_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b110111010;  //node 442
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00001_00010_00000_00010_11110_00001_00010_00001_00001_11111_11110_11111_00011_00001_00001_00000_00010_00000_00000_11111_00000_11111_00000_11111_00000_00001_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b110111011;  //node 443
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00001_00010_00000_00010_11110_00001_00001_11111_00000_00000_00000_00000_00010_00000_00000_00010_00000_00000_11110_00001_00010_11111_00000_11110_00001_11111_00001_11110_11111;

		#2
		WriteAddressSelect <= 10'b110111100;  //node 444
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_11111_00000_00001_00001_00000_00000_00010_00000_00000_00000_11110_00010_00000_00001_00001_11111_11110_00000_00000_11111_11110_00001_11111_11110_11111_00000_11111_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b110111101;  //node 445
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_00000_00010_00001_00001_00001_11111_00000_11110_11111_00001_11110_00001_00001_00000_00001_00001_11111_00011_00011_00000_00000_00001_11111_00000_11111_11111_00000_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b110111110;  //node 446
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00001_11111_00000_11111_00000_00000_11111_11111_00000_00000_00000_00001_00000_00000_00001_00000_11111_00001_00001_00000_00001_11111_00000_00010_11111_00001_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b110111111;  //node 447
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_11111_00001_00000_00001_11111_00000_11111_00001_00001_11111_00001_00001_00001_00000_00001_11111_00001_11111_00001_00001_11111_00001_00000_00001_00001_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b111000000;  //node 448
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00000_00000_00000_00010_00000_00000_00000_00000_11111_00001_00000_00001_00001_11111_11110_00001_00000_11110_00000_00001_00001_00001_00001_00001_00000_00001_00010_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b111000001;  //node 449
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_00000_00000_00001_00000_00001_00000_00000_00010_11111_00001_00000_00000_11111_00000_00000_00000_11111_00000_00010_11111_11111_00000_11111_00000_00000_00000_11110_11110;

		#2
		WriteAddressSelect <= 10'b111000010;  //node 450
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00000_00010_00010_00010_00001_00001_00001_00000_11110_11110_00010_11111_11111_11110_00010_00000_00010_00000_11111_11111_00000_00010_00000_00001_11111_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b111000011;  //node 451
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_00000_11111_11110_11111_00000_00000_00001_11111_11111_00010_11110_00000_00001_00000_11111_00000_11111_00001_11111_11110_00001_00010_00010_00001_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b111000100;  //node 452
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_11110_00000_00000_00001_11110_11110_00001_11111_11110_00000_00000_00001_00001_00000_00000_00000_00010_11111_11110_00000_00000_00001_00010_00000_00011_00000_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b111000101;  //node 453
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00000_00000_00001_00010_00000_00001_00001_11110_00000_11111_00000_00001_00010_00000_00000_00001_00000_00010_11111_11110_00000_00001_00010_00000_11111_00010_00000_11110_11110;

		#2
		WriteAddressSelect <= 10'b111000110;  //node 454
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11111_00010_11111_11111_00001_11111_11101_00010_00000_11111_00000_11110_00000_00001_00001_11111_11110_00000_00110_11110_00001_00001_00000_00000_00000_00000_11110_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b111000111;  //node 455
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_11110_11111_11110_00001_11111_00000_11111_00001_11111_00010_00001_11110_00000_00011_00010_00010_00010_00001_11110_00001_11111_00000_00001_00000_00001_00000_11111_11110_00010_11111;

		#2
		WriteAddressSelect <= 10'b111001000;  //node 456
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00001_11110_00000_00000_00001_11111_00000_00001_00000_00000_11111_00000_00001_00100_00001_00000_00010_00001_11100_00001_00000_11111_11111_00010_00001_00001_00001_11110_00010_00010;

		#2
		WriteAddressSelect <= 10'b111001001;  //node 457
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00010_00000_00001_00001_11111_11110_00000_00000_00010_00000_11111_00010_11111_11111_00010_00001_11110_11111_11010_00001_11110_00000_11110_00001_11111_11110_00000_11110_00010_11111;

		#2
		WriteAddressSelect <= 10'b111001010;  //node 458
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00000_00000_00000_11110_00000_11111_11110_00001_00000_11111_00000_11110_00000_00000_11100_11111_00000_00010_11111_00000_11110_00001_00000_11101_00010_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b111001011;  //node 459
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_00000_00001_00010_00001_00000_00001_11111_11111_00000_00010_11111_00001_11101_00010_11111_11110_00000_00011_11111_00001_11111_00000_00000_11111_11110_00001_00000_00010_11111;

		#2
		WriteAddressSelect <= 10'b111001100;  //node 460
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_11111_00001_00001_00010_00000_00000_11110_11111_00001_00100_11110_00010_11111_00010_00001_00001_11111_00010_11111_00010_11111_00001_11110_00000_11111_11111_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b111001101;  //node 461
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00000_11111_00010_11111_00001_00000_11110_11110_00010_00001_11110_00100_11110_11111_00000_00000_11110_00010_00000_00001_11111_00000_11111_00000_00000_11111_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b111001110;  //node 462
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00001_00001_00011_00010_00010_00000_11110_00010_00001_00010_11110_00000_11111_00000_00000_00010_00001_00000_00001_00000_00010_00010_11110_00001_00000_00000_00000_11110_00001;

		#2
		WriteAddressSelect <= 10'b111001111;  //node 463
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11111_11111_00000_00010_00001_00010_11110_11111_00001_11111_00010_11110_11111_11111_00000_00000_00010_11111_00010_00000_00010_11110_00010_11111_00000_11111_11111_11110_00001_00001;

		#2
		WriteAddressSelect <= 10'b111010000;  //node 464
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_11110_00001_00010_11111_00011_00000_11111_11111_00010_00001_00001_00000_11111_00001_00000_00010_00000_00001_00001_00010_11111_00010_00000_00010_00000_11111_00010_11111_00010;

		#2
		WriteAddressSelect <= 10'b111010001;  //node 465
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_00010_11111_00001_00001_00001_11110_00001_11111_11110_11111_11111_11110_00001_00001_00000_11110_00001_00001_11111_11111_00010_11111_00010_11111_00000_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b111010010;  //node 466
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11111_11111_00000_00000_00000_00010_11110_00001_11110_00001_11101_00001_00010_00000_11111_00000_00001_11111_11111_11111_11110_00001_00001_00001_00001_00000_00001_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b111010011;  //node 467
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_11110_11111_00010_11110_00001_11111_11111_11111_00000_00000_11111_11110_00000_11111_00001_00010_00001_11110_00000_11111_11111_00010_00001_11111_00001_00010_00001_00010_00001_11110;

		#2
		WriteAddressSelect <= 10'b111010100;  //node 468
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00000_11111_00001_00000_00001_00000_00000_00010_11111_11110_00000_11111_00000_00001_11110_00000_11110_00001_00001_11110_00000_00001_00001_00000_11111_00010_00000_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b111010101;  //node 469
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00010_11111_11110_00000_11111_11110_00000_00010_00000_00000_11110_00000_11110_11111_11110_11111_00001_00001_00000_11111_00000_00000_00000_00001_00000_00000_11111_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b111010110;  //node 470
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00011_00001_00000_00001_00000_11111_00011_00001_00001_00000_00000_00000_00000_00011_00010_00000_11111_00010_00000_11110_00000_00010_11111_11111_00001_00010_11110_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b111010111;  //node 471
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11010_00000_00000_00010_00000_00000_11110_00000_00010_11111_11110_00001_00010_00001_00011_00000_11111_00000_00000_00000_11110_11111_00000_00001_00000_11111_00000_11110_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b111011000;  //node 472
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11110_00000_00001_00000_11111_00010_00000_11110_00001_11111_00001_00010_00001_00001_00000_00010_00001_00000_11110_00001_00001_11111_00000_11111_11111_00000_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b111011001;  //node 473
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11111_00000_00001_11111_00001_11111_00001_11111_00010_00001_00000_00001_00000_00010_00000_00000_11111_00001_00000_00000_00000_00001_11111_11111_00000_00000_00000_11110_00010_00001;

		#2
		WriteAddressSelect <= 10'b111011010;  //node 474
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00001_00001_11111_11111_00001_00001_00000_00010_11111_00001_00001_11111_00001_00000_11111_00001_11111_00001_00000_00000_11111_00001_11111_00000_00000_11111_00010_11111;

		#2
		WriteAddressSelect <= 10'b111011011;  //node 475
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00000_11111_00001_11111_00001_11111_00000_00000_11111_00000_11110_00001_00000_00000_11111_00001_00001_11111_00001_00000_00001_00000_00000_11111_00000_00000_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b111011100;  //node 476
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00001_00001_00000_00000_00000_00000_00000_00000_00001_00001_00000_00000_00010_00000_00001_00000_00000_00010_00000_00000_11111_00010_00000_00000_00001_00000_11110_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b111011101;  //node 477
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00001_11111_00000_11111_00000_00001_00001_00000_00000_00001_00000_00001_11111_00000_00010_00010_00000_00000_00001_11111_00000_11111_00000_11111_00001_11111_00001_11110_11111;

		#2
		WriteAddressSelect <= 10'b111011110;  //node 478
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11110_00000_00001_00000_00001_11111_00000_11111_00001_11110_00000_00000_11111_11111_00000_00000_00000_00010_00000_00000_00000_00000_11110_11111_00001_00000_00000_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b111011111;  //node 479
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11110_00001_00010_00001_00000_00001_00000_11110_00000_11111_00000_00000_00010_00001_00001_00001_00000_00000_00001_00000_00000_00000_11110_00000_11111_00001_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b111100000;  //node 480
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_00010_11111_11110_00001_00000_00010_00000_00000_11110_00000_11111_00010_00001_00001_00000_00010_11111_00001_11111_00000_00001_00001_00010_00000_11111_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b111100001;  //node 481
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_11110_00000_00000_00000_11111_11111_00000_00001_11110_11111_11111_00001_00010_00000_00000_00000_11111_00010_11110_11111_00001_00010_00010_00001_11110_11111_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b111100010;  //node 482
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11101_00000_00001_11111_00010_00000_11111_11110_11111_00000_00000_00000_00000_00001_00010_00010_11111_00000_11111_00011_11110_00000_11111_00010_00010_00000_00001_00001_11110_00001_00010;

		#2
		WriteAddressSelect <= 10'b111100011;  //node 483
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00000_11111_00000_00000_00000_00000_00001_11111_00001_00001_00001_11111_00000_00001_00001_00011_00001_11111_00001_00001_00000_00000_00001_00010_00000_00010_00000_00011_00001;

		#2
		WriteAddressSelect <= 10'b111100100;  //node 484
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00001_00000_11110_00001_11111_00000_00000_11110_00010_00000_00001_00010_00001_00010_00010_00000_00000_11100_00010_00000_00001_00000_00010_00000_11111_00000_11110_00001_11111;

		#2
		WriteAddressSelect <= 10'b111100101;  //node 485
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00000_11111_00001_00010_11110_11111_11110_11110_00000_00001_11110_00001_11111_00001_11111_00001_11110_00010_11101_00001_11111_00000_11110_00001_00000_11110_00010_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b111100110;  //node 486
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11111_00000_11111_00001_00000_00000_00000_11110_00001_00000_11110_00010_11111_11110_11111_11111_10111_00000_00000_00010_11110_00001_00000_00011_11111_11110_00010_11111_11110_00000;

		#2
		WriteAddressSelect <= 10'b111100111;  //node 487
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11110_00010_00100_00001_11111_11111_00000_11111_11111_00000_00010_00001_11111_00001_00000_11111_11110_00011_00001_00000_00001_11111_00000_00000_00000_00010_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b111101000;  //node 488
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11110_00000_11111_00011_00001_11111_00001_11111_00000_00001_11111_00001_00010_11111_00001_11111_00010_11110_00010_11110_00001_11111_00001_00000_00000_11111_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b111101001;  //node 489
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_11111_00010_00010_00001_00001_11111_11111_00010_00001_00000_00001_00000_11111_11111_11110_00001_11111_00000_00000_00001_00001_00000_00000_00000_00001_00000_00001_00000_00010;

		#2
		WriteAddressSelect <= 10'b111101010;  //node 490
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00000_00001_00010_00001_00001_00001_11110_00000_00010_00000_11110_11111_11110_11111_00001_00010_00001_00001_00001_00010_00000_00010_00001_00001_11111_11111_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b111101011;  //node 491
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_11110_00010_00010_11111_00010_00000_11110_00001_00001_11110_11110_00000_11110_00000_11111_00000_00001_00001_00001_00001_00001_00010_00001_00010_00000_00000_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b111101100;  //node 492
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00000_00000_00010_11111_00000_00011_00001_11110_11111_00010_11011_11111_11111_11111_11111_00001_00001_11111_11111_00000_00000_00001_00010_00000_11111_11111_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b111101101;  //node 493
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00000_11101_00010_11110_00000_00000_11111_11111_11110_00001_11110_11111_00000_00000_11110_00000_00001_11110_00001_11111_00000_00000_00010_00001_00001_00000_00001_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b111101110;  //node 494
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_11111_11110_00001_11101_11111_00000_11111_00001_11111_00010_00000_11110_00010_00000_11111_00010_11111_00000_00000_00000_00001_00010_00001_00001_00010_11110_00000_00010_00000_11110;

		#2
		WriteAddressSelect <= 10'b111101111;  //node 495
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_11111_00000_11101_00001_11111_11111_11111_00001_11110_11111_00000_11110_00001_11111_11111_00000_11110_11111_11111_00001_00010_00000_00000_11111_00000_11110_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b111110000;  //node 496
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11111_11111_00001_11111_00010_00000_00000_00001_00001_11111_00010_00001_00010_00001_00000_00000_00001_00000_00000_00000_00011_00001_00001_11110_11110_00011_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b111110001;  //node 497
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_11111_11111_00000_11111_11111_00000_11111_00001_00000_11111_00000_00001_00010_00000_00010_00010_11111_11110_11110_00001_00001_00010_00000_00001_11111_00000_00001_11110;

		#2
		WriteAddressSelect <= 10'b111110010;  //node 498
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11111_00000_00000_00001_11111_00000_00001_00001_00001_00000_00000_00001_00001_00001_00000_00001_00000_00000_11111_00000_00001_11111_11111_11111_00000_11111_00001_11110_11110;

		#2
		WriteAddressSelect <= 10'b111110011;  //node 499
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11011_11111_00000_00000_00010_00001_11111_00010_00010_00000_00000_00001_00001_00000_00010_00000_11111_11111_00000_11111_11111_00001_00001_00001_00001_00001_00001_11111_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b111110100;  //node 500
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11010_00000_00000_11111_00010_00000_00000_00001_00000_00010_00000_11111_11110_00000_11111_00001_00001_11111_11111_00001_00001_00001_00010_00010_11110_00000_00000_00000_00000_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b111110101;  //node 501
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00000_00000_00001_11111_00000_11111_11111_00000_00001_00001_00001_00000_00001_00000_11111_11110_00010_00000_00010_00001_11111_00000_00001_11111_11110_00001_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b111110110;  //node 502
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_00001_11111_11111_00000_11111_00000_11110_00010_00000_11111_00000_11111_00001_00000_00000_00000_00000_00010_00001_00001_00000_00000_11111_11111_00010_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b111110111;  //node 503
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_11111_00001_00001_00000_11111_00001_11111_00000_00000_00000_00010_00000_00001_00000_00010_00000_00001_11111_00000_11111_00000_00001_00001_00000_00001_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b111111000;  //node 504
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_00000_00001_00000_11110_00001_11110_00000_00001_00000_11111_11111_00000_00000_00001_00001_00000_00001_11110_00000_11111_00001_00000_00001_11111_11111_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b111111001;  //node 505
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_11111_00000_00000_00001_00001_00001_00000_00000_11111_00001_00000_00000_00001_11110_11111_00000_00001_11111_00000_00000_11111_00000_00001_11110_00000_00000_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b111111010;  //node 506
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_11111_00000_00001_00001_00000_00000_00000_00001_00001_00001_11111_00000_00000_00000_00000_00001_00001_00001_00001_00001_00010_00010_00000_00000_11111_11111_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b111111011;  //node 507
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00010_00000_00001_00000_00001_00000_00001_00000_00000_00001_11111_00010_11111_00001_11111_00000_00010_00000_11110_00000_00000_11110_11111_00000_00001_11111_00010_00000_11110_00010;

		#2
		WriteAddressSelect <= 10'b111111100;  //node 508
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11110_00000_00001_00001_00001_00000_11110_00001_11111_00000_00000_00000_00001_00010_00000_00000_11110_00001_00010_11111_00000_00000_00001_00000_00000_00010_00001_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b111111101;  //node 509
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_11111_00010_00001_11111_00000_00000_00001_00010_11111_00000_00010_11111_00010_00010_00010_11111_00000_00000_00010_11110_11111_00001_00001_00010_00000_00010_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b111111110;  //node 510
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_00000_11111_00001_00000_11111_11111_00000_00001_00000_00001_11111_00000_00010_00010_00001_00001_00001_00010_11111_00000_00000_00001_00011_00001_00000_00001_11110_00011_00001;

		#2
		WriteAddressSelect <= 10'b111111111;  //node 511
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00001_00001_00010_00000_00000_00010_00010_00001_00001_00001_00000_00001_00011_00010_00001_00011_00010_11110_11111_00001_00001_00000_00010_00000_00010_00000_00000_00010_00010;

		#2
		WriteAddressSelect <= 10'b1000000000;  //node 512
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_11111_00001_11111_00001_00001_00001_00010_00010_00000_00001_00000_00000_11111_00001_11111_00000_00000_00010_11110_00000_00010_00000_00000_00011_11110_11110_00000_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b1000000001;  //node 513
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_11111_00000_00000_11101_11111_11110_00000_00000_00001_11111_00010_00001_00001_00001_11111_11110_00001_11100_00011_00001_00001_00000_00011_11111_00000_00001_11110_00001_00000;

		#2
		WriteAddressSelect <= 10'b1000000010;  //node 514
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_11110_00001_00000_11111_11111_00001_11111_11111_11111_11111_11110_00001_00000_00000_00001_10101_00010_00000_00010_00000_00000_11111_00011_00000_11110_00001_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1000000011;  //node 515
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_11111_11111_00000_00000_00000_11110_00001_00000_00000_00010_11111_00000_00010_00001_00001_11110_11110_00000_00010_11111_11111_00000_11111_00011_11111_00000_00010_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1000000100;  //node 516
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_11111_00001_00010_00000_11111_00001_11111_11111_00000_00000_11111_11111_00000_11111_00000_00010_11111_00011_11110_00000_00001_11111_00001_00000_11111_00001_11110_11111_00010;

		#2
		WriteAddressSelect <= 10'b1000000101;  //node 517
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00000_11111_00000_00001_00001_00001_11111_00000_00001_11110_00010_00000_11110_00000_00000_00010_11110_11111_00001_00010_00000_00001_00001_00010_11110_00000_00000_00001_00010;

		#2
		WriteAddressSelect <= 10'b1000000110;  //node 518
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11111_11111_00001_00010_00000_00001_00010_00000_00000_00001_00000_11110_00000_11111_00001_00001_00001_00000_00001_11111_00000_11111_00010_00000_00001_11111_11111_11110_00010_00001;

		#2
		WriteAddressSelect <= 10'b1000000111;  //node 519
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00010_00001_00010_00000_11110_00001_00000_11111_00001_00010_11110_00001_11110_11110_00000_00000_00001_00000_00001_00000_00010_00000_00000_00001_00010_00001_00001_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1000001000;  //node 520
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_11110_00010_11110_00000_00001_11110_00000_00001_00001_11110_11111_00001_11110_11111_00001_11111_11111_00000_11111_00000_11111_00000_00000_00001_11110_00001_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1000001001;  //node 521
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_11111_00010_11110_11111_11111_00000_00010_11111_00000_00000_11111_00010_11110_00000_00000_00001_11111_00010_00001_00000_00000_00001_11111_00001_00001_00000_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b1000001010;  //node 522
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_00010_11111_11111_11110_00000_11111_00001_00000_00000_11110_00010_11111_11111_00000_00000_00000_00000_11111_00000_11111_11110_00010_00000_00001_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1000001011;  //node 523
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00010_00000_00000_11110_00010_00001_00000_00000_11111_11111_11111_00000_00000_11111_00000_11111_00001_00000_00001_11110_00001_00001_00010_11111_00000_00000_00001_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b1000001100;  //node 524
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00001_11111_00000_11111_00000_11111_00001_00000_00000_11111_00000_00001_00001_00000_00000_11111_00000_00000_00000_00000_11111_00001_00001_00001_00010_00010_11111_11110_11111_00000;

		#2
		WriteAddressSelect <= 10'b1000001101;  //node 525
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11110_00000_11110_00010_00001_00001_00001_11111_11111_00001_11111_00001_00010_00010_11111_00000_00000_11111_00000_00000_00000_00001_00000_11110_00100_11110_11110_11111_11110;

		#2
		WriteAddressSelect <= 10'b1000001110;  //node 526
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_00000_11111_11111_00001_11111_00000_00010_11111_00000_00000_00000_00000_00011_00000_11111_11111_00001_00000_00000_00000_00001_00000_00000_11111_00001_11101_11110_11111_11111;

		#2
		WriteAddressSelect <= 10'b1000001111;  //node 527
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11011_00001_00010_11110_00001_00000_11111_00001_00010_11111_11111_00001_00010_00000_00000_11111_00001_11111_00001_00000_11111_00000_00000_00001_11111_00000_11110_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1000010000;  //node 528
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_11110_00001_11110_00001_00001_11111_00001_00000_11111_00000_00000_00000_00010_00000_11110_11111_00001_00000_11111_00000_00010_00010_11111_00000_00001_00000_00001_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000010001;  //node 529
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_11111_00000_11111_11111_00001_00000_00001_00010_00000_00010_00000_00000_00001_00000_11111_00000_00001_00000_11111_11111_11111_00000_11110_00001_00010_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b1000010010;  //node 530
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_00001_11110_00001_11111_11111_00001_11110_00001_00010_00000_11111_00001_11111_00001_11111_11111_00000_11111_00001_00000_11111_00000_00001_11111_00000_00000_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1000010011;  //node 531
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00000_11111_00001_11110_00001_00000_00000_00000_00000_00001_11111_11111_00000_11110_11111_00010_00000_00000_00001_11111_00000_00001_11111_00000_00001_11111_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1000010100;  //node 532
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00001_00001_00000_00001_11111_11111_11110_11111_00000_11110_11111_11111_00000_00000_00000_11110_00001_00000_11111_11111_00000_00001_00000_00010_00001_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1000010101;  //node 533
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_00000_00000_00000_00001_00000_00000_00000_00000_00001_11111_00001_11111_00000_11111_00001_00000_11111_11111_00001_00001_00000_00001_00001_00001_11111_11110_00001_11110_11111_11111;

		#2
		WriteAddressSelect <= 10'b1000010110;  //node 534
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00001_11111_00000_00001_00000_00001_00000_00001_00000_00000_00000_11111_11111_11111_00000_11110_00000_00000_11111_11111_11111_11110_00001_00000_00000_00000_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1000010111;  //node 535
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00010_00000_00000_11111_11110_00001_00000_00001_00001_00001_00001_00000_00000_00001_00001_00000_11111_00001_00000_00000_00001_00001_11111_00001_00001_00000_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1000011000;  //node 536
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00010_00001_00000_00001_00000_11111_11111_00001_11110_11111_11111_00010_00001_00001_00000_00000_00001_00010_00001_00011_11111_11111_00000_00000_00010_00000_00001_11110_11111;

		#2
		WriteAddressSelect <= 10'b1000011001;  //node 537
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_11111_00000_00010_00001_00000_11111_00000_11111_11111_11111_00000_00001_00001_11111_00010_00001_00010_11101_00000_00001_00001_00010_00001_00000_00000_11111_11110_00000;

		#2
		WriteAddressSelect <= 10'b1000011010;  //node 538
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00001_00000_11110_00001_00000_11111_00000_00001_00001_00000_00001_00000_00001_00010_00001_00001_00010_00010_11101_00000_00001_00001_00011_00000_00010_00001_00001_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000011011;  //node 539
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00010_00001_00001_00010_00000_00001_00000_00001_00010_00001_11110_00001_00001_00011_00010_00001_00100_00010_00000_11111_00000_00000_00000_00101_11111_00000_00000_11110_11111_00001;

		#2
		WriteAddressSelect <= 10'b1000011100;  //node 540
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_11110_00010_00000_11111_00000_11111_11110_00000_11111_00000_11111_00001_11111_00000_00010_00010_11110_00010_00000_00010_00000_00001_00000_00001_11111_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1000011101;  //node 541
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11110_11111_00000_00001_00000_00001_11110_00000_00001_11110_00001_11111_00000_00000_11111_11111_00000_11110_00010_11111_00001_00001_00011_11110_00000_00001_11111_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000011110;  //node 542
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_11110_00001_00010_00001_11111_11110_00000_11110_00010_00001_11110_11111_00001_00000_00000_00000_11001_00000_11111_00001_00001_11111_00001_00010_00000_11110_00010_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b1000011111;  //node 543
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_11110_00001_11110_00000_11111_00001_11110_00001_00010_11110_00000_00010_00010_00000_00000_10110_11111_00010_00010_11111_11110_00001_00000_00001_11111_00000_11110_00000_11111;

		#2
		WriteAddressSelect <= 10'b1000100000;  //node 544
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_11111_00010_00001_00001_00000_00000_00000_11110_11110_00001_00000_00000_00001_11110_11110_11110_11110_00010_00000_11111_00010_00001_11111_11111_00000_00000_11111_00001_11110;

		#2
		WriteAddressSelect <= 10'b1000100001;  //node 545
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_11111_00000_00000_00000_11111_00001_00000_00001_00000_11110_00000_11110_11111_00000_11111_00001_00000_00000_00000_00000_11111_00001_11111_00000_11110_11110_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1000100010;  //node 546
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_00001_00001_11111_11111_00000_11110_00001_00001_11111_11111_11110_11110_00010_00001_00000_00000_00000_11111_00010_00010_00000_11111_00000_00000_11111_00000_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000100011;  //node 547
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00010_00000_00010_11110_00001_11110_11111_00001_11111_00001_11100_11111_11110_11111_11110_00000_00000_11111_00001_11111_00000_00010_00010_00000_00001_11110_11110_11110_00000_11111;

		#2
		WriteAddressSelect <= 10'b1000100100;  //node 548
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_11110_00010_11101_11111_11111_00001_11111_00000_00001_11110_00001_00000_11110_11111_00000_00000_00001_00001_11111_00001_00000_11110_00001_00001_00000_11111_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b1000100101;  //node 549
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_00001_00001_11111_00000_00000_00010_00001_11111_11110_11111_00000_00010_11111_11111_00010_11110_11111_00000_00000_00001_00011_00000_00000_11110_11111_00000_00000_11110_11110;

		#2
		WriteAddressSelect <= 10'b1000100110;  //node 550
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_00001_11111_00010_11111_00010_00000_00001_00001_11111_00000_11111_00000_00001_00010_00000_11111_00001_00001_11111_00001_11111_00001_11110_00010_00000_00000_11111_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1000100111;  //node 551
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11101_00000_00010_11111_00001_11110_00000_11110_11111_11111_00001_11111_00000_11111_00001_11111_11110_00000_11111_00010_00001_00000_00000_00010_11111_00000_11110_00001_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1000101000;  //node 552
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_00000_00000_11111_11111_00000_00000_00001_00001_11111_00001_11110_00010_00001_00000_00000_00001_11111_11111_11110_00001_00000_11111_00000_00000_00010_11110_11110_11111_11111;

		#2
		WriteAddressSelect <= 10'b1000101001;  //node 553
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_00000_00000_00010_00000_11110_00000_00000_00000_00000_00001_00001_00000_00010_00000_00000_11111_00010_11111_11111_00001_00010_00001_11111_11111_00001_11110_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b1000101010;  //node 554
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00000_00000_00000_11110_11101_00001_00001_00010_00000_00001_00000_00001_00010_11111_00010_00001_00001_11111_11111_00001_00000_00001_11111_00000_00000_00000_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b1000101011;  //node 555
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00001_00000_11111_00001_00000_11111_11111_00000_00000_11111_11111_00000_00000_11111_00001_00000_00001_00001_00000_11110_11111_00000_00010_00000_11111_00000_11111_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b1000101100;  //node 556
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11101_00001_00000_00000_00000_00000_00000_00001_00000_00000_11111_00001_00001_11111_00010_00001_11111_00000_11111_11111_00001_11111_00010_00000_00000_11111_00000_11111_00000_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000101101;  //node 557
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_11111_11111_00001_00000_00000_00000_00001_11111_00000_11111_00000_00000_11111_00000_11111_00000_00001_00000_00000_00001_00001_11110_11111_00000_00000_11111_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b1000101110;  //node 558
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_11111_00001_00000_11111_00000_00000_00010_00000_11110_00000_00000_00001_00000_00000_11111_11110_11111_11111_00000_00000_11111_00001_11111_11111_00001_00010_11111_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1000101111;  //node 559
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00001_00000_00000_11111_00000_00001_00001_11111_00000_11111_00001_11111_00010_00010_00000_00001_11111_11111_00001_00001_00001_00001_00000_00000_00001_11111_00000_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1000110000;  //node 560
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_00001_11110_00001_00000_11111_00000_00000_00001_00001_00000_00000_00001_00000_00000_00000_11111_11110_00001_00000_00010_11111_11111_11111_00001_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1000110001;  //node 561
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00001_00001_11110_11111_00001_00000_00000_00010_11111_00000_11111_00001_00001_00000_00000_00000_00000_11111_11111_00000_11110_11111_00001_00010_00001_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1000110010;  //node 562
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11111_00000_00010_00000_00000_11111_00001_00001_00000_00001_00000_11111_00000_00001_00000_00000_00000_00000_11110_00000_00000_00001_00000_11111_00000_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1000110011;  //node 563
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_00001_11111_11110_00010_11110_00001_00001_11111_11110_11111_11110_11111_11110_00000_00001_00000_00000_00000_00001_11110_11111_00000_11110_00000_00000_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1000110100;  //node 564
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00010_00001_00000_00000_00000_00000_00000_00000_11111_00000_00000_00000_11111_00001_11111_00001_00000_00010_00001_00001_11111_00001_00010_11111_11101_11111_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1000110101;  //node 565
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_00000_11111_11111_00000_00000_00000_11111_00001_00000_00010_00101_11111_11111_00000_00010_00000_00000_11111_00001_00000_00010_11111_00001_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1000110110;  //node 566
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00001_00000_00001_00001_00000_00001_00010_00001_00001_00000_11111_11111_00000_00000_00001_00010_00010_00001_11111_11110_00001_00000_00001_11110_11110_00000_11111_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000110111;  //node 567
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_00001_00010_00000_00001_11111_00001_11111_00001_00000_00000_00000_11110_00001_00010_00001_00001_00101_00010_11101_00001_00001_00001_11111_00010_11111_00001_00001_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b1000111000;  //node 568
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00001_11111_11110_11110_11111_11111_00001_00001_00000_11110_00010_11110_00001_00000_00010_00001_00010_11110_00010_00000_11111_00010_00010_00000_11111_00000_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b1000111001;  //node 569
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_00000_00000_00000_00000_11111_00011_00000_11111_00001_11110_00000_00010_11111_11111_11111_00000_00001_11011_00001_00010_00000_00010_00010_11111_11110_00000_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b1000111010;  //node 570
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_00000_11111_00001_00001_00010_00000_00001_00001_11111_00010_00000_00001_11111_11110_11011_00000_00000_00001_00010_00001_11111_00010_11111_11111_00010_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1000111011;  //node 571
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_11111_00001_11110_00000_11111_00000_00000_11111_00010_11110_11111_00001_11111_00001_00000_11111_11011_11111_11110_00001_11111_00000_00010_11110_11101_00000_00001_00010_00001;

		#2
		WriteAddressSelect <= 10'b1000111100;  //node 572
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_11110_00001_11111_11110_00000_11111_00001_00000_11111_11111_00000_00000_00010_00000_11111_11111_00010_11110_00001_00000_00001_00001_00000_11111_00000_00001_00010_11111;

		#2
		WriteAddressSelect <= 10'b1000111101;  //node 573
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00010_00000_00001_11110_11111_00001_00001_11111_00001_00001_00001_00000_11111_00001_00000_11110_00000_11111_00010_11101_00000_00001_00010_11111_00011_00001_11110_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b1000111110;  //node 574
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00010_00001_00001_11110_11110_00000_00001_00001_00001_00010_00000_00000_11111_11110_00000_00000_00000_11111_11111_11110_00000_00001_00000_11111_00000_00000_00000_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b1000111111;  //node 575
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00000_11111_00001_00000_00001_11110_00001_00001_11101_00001_00001_11110_11111_00000_00000_11110_00010_00000_00000_11110_00010_00001_00000_00001_00000_00001_00000_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b1001000000;  //node 576
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00010_11111_00000_11111_11110_00000_00001_00010_11110_00001_11111_00001_00000_11110_00000_00001_00000_11110_00001_11111_00001_00010_11111_00000_00000_11111_11111_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001000001;  //node 577
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00001_00000_00010_11110_00001_00000_00001_00001_00001_00001_11111_00001_11111_11110_00000_00000_00010_11111_00001_00000_00000_00000_00000_11111_11111_00000_11110_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b1001000010;  //node 578
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00001_00001_00001_11111_00000_11111_00000_11110_11111_00001_11110_11111_00010_11111_11111_00001_00010_00000_11111_11111_00001_00000_00001_00000_00001_00000_11110_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1001000011;  //node 579
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_11111_11111_11110_00000_00001_00010_00011_00000_00000_00001_11111_11111_00001_00001_00000_00000_00010_00000_11110_00000_00000_00001_11111_00000_00001_11110_11110_00010_11110;

		#2
		WriteAddressSelect <= 10'b1001000100;  //node 580
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11101_00000_00010_00000_00001_00000_00010_00001_11111_11111_00010_11111_00000_00000_00000_00001_00000_00001_00000_00000_00000_00000_11111_00001_00000_00000_11111_00001_11110_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001000101;  //node 581
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00010_11111_00000_00001_00000_00010_11111_00001_00000_11110_11111_11110_00010_00010_00000_11111_11110_00010_11111_00000_00000_00010_11111_00000_11111_00010_11110_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b1001000110;  //node 582
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11101_00001_00000_00010_00001_00000_00001_00000_11111_00000_00000_00000_00000_11111_00000_00000_00001_00001_00000_00001_00000_00000_11111_00001_00000_11111_00000_00010_11111_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1001000111;  //node 583
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_11111_11111_11111_00001_11111_00010_00001_00000_00000_00000_00000_00010_00001_11110_00001_00010_11111_00001_11110_00001_00000_11111_00010_00001_11110_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1001001000;  //node 584
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11111_11111_00000_00000_00001_00000_11111_00010_00001_11111_00000_00000_00000_00001_11110_00001_11110_11111_00000_11111_00001_00001_00010_00000_11111_00010_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b1001001001;  //node 585
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11110_00000_00010_11111_00001_11111_11111_00000_11111_11111_11110_11111_00001_00000_11110_11110_00000_11111_11110_11111_11110_00000_11110_00000_00010_00010_00001_11110_00001_11110;

		#2
		WriteAddressSelect <= 10'b1001001010;  //node 586
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00001_00001_00000_00000_00000_00001_00001_11111_00000_00010_11111_00001_11110_00001_11111_00000_00001_00001_11111_00000_11111_11111_00000_00001_00000_11111_00001_00001_00010;

		#2
		WriteAddressSelect <= 10'b1001001011;  //node 587
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_00001_00010_11111_00001_00001_11111_00001_00010_00000_00000_00000_00000_00000_00010_11111_00001_00000_00000_11111_11111_00000_11111_00010_00000_11111_00000_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b1001001100;  //node 588
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11110_11111_00010_00000_00000_00000_11111_00000_00010_00000_00000_00000_11111_00010_00000_00001_00000_11110_11111_00001_11111_11111_00010_00000_00001_00000_00010_11111_00001;

		#2
		WriteAddressSelect <= 10'b1001001101;  //node 589
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_11111_11111_11111_00001_00000_11110_00010_00001_00000_00001_00000_00000_00000_11110_00010_00000_00001_00000_00000_00001_11111_00010_00001_11111_11111_00000_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b1001001110;  //node 590
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11110_00000_11111_00000_00001_11111_00001_11111_11111_00000_00000_11111_00001_00000_11111_00001_00010_00001_00001_11110_00010_00001_00001_11111_00001_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001001111;  //node 591
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11110_00010_00001_11110_00010_00001_11111_00000_00001_11111_00010_00000_00000_00000_00000_11111_00001_00001_00001_00001_11111_00000_00000_11111_00001_11111_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001010000;  //node 592
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11101_11111_00000_00001_00001_00001_00000_11111_00000_00000_00001_00000_11110_11110_11110_00000_11111_00001_00001_00001_11110_00001_00001_11111_00000_00000_11111_00010_00001_11110_00001;

		#2
		WriteAddressSelect <= 10'b1001010001;  //node 593
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00000_11111_11110_11111_00000_00001_00001_00001_11110_00010_11111_00001_00010_00010_11111_00001_00010_11111_11110_00000_00001_00000_00001_00000_00000_00000_00010_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001010010;  //node 594
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_11110_00001_00000_00000_00001_11111_00000_00010_11110_00010_11111_00010_11110_00000_00000_00001_00001_00001_00001_00000_11111_00001_00001_00001_00000_00001_00000_11011_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001010011;  //node 595
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11110_00001_00010_11111_00000_00001_11111_00000_11111_00000_11111_00001_11110_11111_00000_11110_00010_00010_11111_00001_00000_00000_00010_00010_11111_00000_00010_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1001010100;  //node 596
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_00000_00000_11111_00001_00000_00001_00000_00001_00010_11111_00000_00000_00001_11111_00001_00000_00001_11111_00010_11110_00010_00000_00010_00000_00000_00010_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001010101;  //node 597
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_00000_00000_00000_00001_11111_00000_00000_00010_11111_11110_00001_00001_00000_11111_11110_11110_00000_11110_00010_00001_00000_00001_00000_11111_00001_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001010110;  //node 598
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_00001_00001_00001_11110_11110_11111_00000_00001_11110_00010_11110_11111_00000_11111_11100_11111_11111_00010_00010_11110_00000_00000_11111_11110_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001010111;  //node 599
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_00001_11110_00000_00001_00000_11111_00000_11111_11110_11111_00000_00000_00000_00001_11110_11111_00000_00010_11110_00001_00000_11111_11110_00010_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1001011000;  //node 600
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_00000_00001_11111_11110_00010_11110_00000_00000_11111_00000_11110_00000_00001_00000_00000_11110_00010_11110_00000_00001_00000_00000_11111_00000_11111_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b1001011001;  //node 601
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00000_00001_11111_11110_00001_00010_11111_11111_00000_11110_11110_11111_11111_11111_00000_11111_11111_11101_00000_00001_00000_00000_00001_11111_11111_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001011010;  //node 602
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_00000_00000_00001_11111_00001_00000_00010_00001_00001_00001_00000_11110_11110_11110_00001_00010_00000_11110_11111_11110_00000_11110_00001_00000_00000_00000_00000_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1001011011;  //node 603
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_11110_00000_00000_00000_11110_00001_00001_00000_00010_00000_00000_00000_11110_00001_11111_11111_11111_00000_00001_00001_00000_00000_00000_11111_00001_00000_00000_11110_11110;

		#2
		WriteAddressSelect <= 10'b1001011100;  //node 604
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11101_00010_00000_11110_00010_11110_11111_00000_00000_00001_00010_00001_00000_00001_00000_00000_00001_00001_00001_11111_11111_11110_00000_00000_11111_00010_00000_00001_11111_00001_11110_00010;

		#2
		WriteAddressSelect <= 10'b1001011101;  //node 605
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00001_00000_00001_11111_00000_11111_11111_00001_00000_11111_11110_00001_00010_11101_11110_11111_11111_00000_11111_11110_11111_00000_00000_11111_00001_00000_11111_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001011110;  //node 606
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_00001_11110_00001_11111_00000_00000_00000_00001_00000_00000_00000_11111_00001_00000_11111_00001_11111_00001_00000_00001_00000_00001_00000_00001_11110_00000_11110_00001;

		#2
		WriteAddressSelect <= 10'b1001011111;  //node 607
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_00000_00010_11111_11110_00001_11111_00000_00000_00001_11111_00000_00000_00010_00001_00001_11111_00001_11111_00000_00001_00001_00010_00000_00001_00000_00001_11110_00000_11110_00010;

		#2
		WriteAddressSelect <= 10'b1001100000;  //node 608
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_00001_00001_00000_00000_00000_11110_11111_00000_00010_11110_00000_00000_00001_00010_00010_11111_00000_00001_00000_00010_11111_00001_00000_00000_11111_00010_00000_11110_00001_00010;

		#2
		WriteAddressSelect <= 10'b1001100001;  //node 609
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_00000_11110_00000_11111_11111_00001_00001_11111_00001_11110_00000_00000_11111_00000_00000_00000_00001_00000_11111_00000_00001_11111_00001_11111_11110_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001100010;  //node 610
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_00001_00000_11111_11111_11111_11111_00000_11111_00000_11111_00001_00000_00010_00000_00001_00010_11111_11110_11110_00001_00010_00000_11111_00000_00000_11111_00001_00000;

		#2
		WriteAddressSelect <= 10'b1001100011;  //node 611
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00001_11110_00010_00000_11111_11111_11111_00001_00000_11111_11111_00000_00001_00001_11110_11111_11111_00010_11111_00000_00001_00001_00000_00001_11111_00000_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001100100;  //node 612
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_11110_00000_00001_11111_00001_00000_00000_00000_00000_11111_00000_00000_00001_00000_11111_11111_00000_00010_11111_00000_00010_00001_00000_11111_00000_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001100101;  //node 613
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_11110_00000_11111_11111_00001_00000_11111_00001_00001_00001_11111_00001_00000_00000_11111_00000_11110_00000_00000_11111_11111_11111_11110_11111_11111_00000_11110_00001_11111;

		#2
		WriteAddressSelect <= 10'b1001100110;  //node 614
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00010_00000_00000_00001_00000_11111_11111_00001_00000_11110_00001_11111_00000_00000_11111_00001_00001_11111_00010_00001_11111_11111_00001_00001_11111_00001_00001_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1001100111;  //node 615
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11110_00001_00000_00000_00000_00000_11111_11111_00000_11111_00000_11111_11110_11111_11111_00001_11111_11111_00001_11110_11110_00000_00000_00000_11111_11111_00000_00000_00001_00001_11110;

		#2
		WriteAddressSelect <= 10'b1001101000;  //node 616
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_11111_00000_11111_00010_11111_00000_00000_00000_00000_00000_00000_00001_00000_00001_00000_00000_00010_00000_11111_00000_00000_00010_00001_11111_00001_11111_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1001101001;  //node 617
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00000_11110_00001_00000_00000_11111_00001_00000_11110_00001_11111_11110_00000_11111_11111_00001_00010_00001_00000_11110_00000_00000_11111_00001_00000_11111_11110_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b1001101010;  //node 618
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_00000_00001_00000_00000_00000_00001_00000_00000_00010_00000_00000_00000_11110_00001_11111_00010_00000_00000_00000_11111_11111_11111_00000_00001_11111_00001_00010_11110_00000;

		#2
		WriteAddressSelect <= 10'b1001101011;  //node 619
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_11111_00000_00000_00000_00000_00010_00000_11111_00000_00001_00000_00001_00000_11111_11110_00001_11111_00000_00000_00001_00000_11111_00001_11111_00000_00010_00001_00001;

		#2
		WriteAddressSelect <= 10'b1001101100;  //node 620
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_11111_00010_00000_00000_00001_00010_00001_11111_00000_00000_11111_11110_00001_00001_00001_00010_00000_00001_00001_11111_00010_00001_00000_11111_00000_00000_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b1001101101;  //node 621
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_00000_00000_11111_00001_00000_00001_00001_00000_00000_11111_11111_00000_11111_00000_00010_00001_11110_11111_11111_00001_00001_00000_11111_11111_00000_00000_11110_00010;

		#2
		WriteAddressSelect <= 10'b1001101110;  //node 622
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00000_00010_00010_00000_00000_11111_00010_00001_00001_00000_00000_00000_00000_11111_00000_00000_00000_00001_00000_00001_00000_11111_00001_00010_00000_00001_11110_00000_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b1001101111;  //node 623
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_00001_00001_00000_00000_00001_00000_00000_11111_00000_00001_00001_00010_00000_00001_00000_00001_11111_00010_00000_11111_00010_00001_00001_11111_00000_11110_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001110000;  //node 624
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_11111_00001_00001_00001_00000_00001_11111_00000_11110_00001_11111_00010_00000_00010_00000_00000_11110_00000_11110_00010_00010_00010_00010_00000_00000_00000_00000_00000_00000_00010;

		#2
		WriteAddressSelect <= 10'b1001110001;  //node 625
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00000_11111_00000_00000_11111_11110_00001_00000_00010_11110_00001_00001_00001_11111_00001_00001_00010_11101_00001_00010_00001_11111_00001_11110_00000_00010_00000_11111_11110;

		#2
		WriteAddressSelect <= 10'b1001110010;  //node 626
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_11110_11111_00000_11110_11111_00000_11110_00010_00000_00000_00010_00000_00000_00000_11111_11110_11111_11110_00001_00000_11111_00001_00010_00000_00000_00001_00001_00010_11111;

		#2
		WriteAddressSelect <= 10'b1001110011;  //node 627
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11110_11110_11111_00000_11111_00001_00000_00000_00001_11111_00000_11101_00000_00001_00000_11010_11100_00000_00000_00000_11110_00001_00010_11111_11111_00010_00000_00010_00001;

		#2
		WriteAddressSelect <= 10'b1001110100;  //node 628
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00001_00010_00001_11111_00000_00001_11110_11111_00001_00001_11111_11110_11111_11111_11110_11111_11110_00000_11101_00001_11110_11111_11111_00000_00000_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1001110101;  //node 629
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00001_11111_00010_11111_00000_00011_00000_00000_11111_00000_11110_00000_11110_00000_00001_11110_11111_00000_00000_00001_11110_00000_00001_00001_00000_00000_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1001110110;  //node 630
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_11110_00001_11111_11110_11111_00010_00000_11111_11111_11111_11111_11110_00010_00000_00001_00000_00000_00000_11110_00001_00000_00000_11111_00000_11111_11110_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1001110111;  //node 631
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00010_11111_00001_11111_11111_00010_00000_11111_11111_11111_00000_11110_11111_00001_00000_11110_00000_11110_00000_00001_11110_11111_00000_11111_11111_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1001111000;  //node 632
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_11111_00000_00000_00000_00000_00001_00010_11111_00000_00001_11111_11111_00000_11110_00000_00000_00000_00001_00000_00000_00001_00000_00001_11110_00000_11110_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1001111001;  //node 633
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00000_11111_11111_00001_11110_00010_00001_00000_00000_11110_00001_00000_00000_00000_00001_11111_00000_11111_00000_11111_00001_11110_00001_11110_11111_11111_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b1001111010;  //node 634
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00001_11111_11110_00000_00001_00000_11111_00001_00010_00000_00000_00000_00001_00000_00001_00000_00000_00000_00001_00000_00000_00000_00000_00000_11111_00001_11110_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b1001111011;  //node 635
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11110_11111_11110_00000_00000_11111_11110_00001_00000_00000_11111_00000_00000_00001_00000_11110_00000_00010_11111_00000_00000_00001_00000_00000_00000_11111_00000_11111_11110_00001;

		#2
		WriteAddressSelect <= 10'b1001111100;  //node 636
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_11111_11111_00000_00010_11111_11111_00001_00000_00000_00001_00001_00001_11111_00000_11111_00001_00000_00000_11110_00001_00001_11111_00000_00001_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1001111101;  //node 637
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_00001_11111_00000_11111_00001_00001_00000_11110_11111_00001_00010_00001_00001_11111_00001_00000_00001_11111_00000_00000_00010_00001_11111_00000_00001_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1001111110;  //node 638
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_11111_00000_00000_11111_11111_11110_00001_00000_00000_11111_11111_00000_00000_00000_11111_00000_00010_00000_00001_00000_11111_11111_11111_00001_00000_00000_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b1001111111;  //node 639
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11110_00000_00000_11110_00000_00001_00000_00000_00000_00000_00001_00001_00001_00000_00000_00001_00000_11110_00000_11111_11111_11111_00001_00010_00000_00000_00001_11110_00001_00001;

		#2
		WriteAddressSelect <= 10'b1010000000;  //node 640
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00010_00000_00000_00000_00000_11111_00000_00001_00000_00010_00001_00000_11111_00001_00000_11110_11110_00000_11111_00000_00000_00000_11111_00000_00010_00001_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1010000001;  //node 641
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_11111_11111_00010_00001_11110_00000_00000_11111_00000_11110_11111_00000_00000_00001_11111_00001_00000_00000_00010_00000_00001_00000_00000_00000_00001_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1010000010;  //node 642
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_11111_11111_00001_00000_00000_00001_00001_00000_00000_00001_11111_00001_00001_11111_00001_11111_00001_11111_00000_00000_00001_11110_11111_00000_00001_11111_00001_00000_00001_11110;

		#2
		WriteAddressSelect <= 10'b1010000011;  //node 643
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00000_00000_00000_00001_00000_00010_00000_11111_11111_00000_11111_11110_00000_00000_00001_00000_11111_11110_11111_00010_00001_11111_11111_11111_00000_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010000100;  //node 644
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_00001_00000_00000_00001_00000_11111_00000_00010_00001_11111_00001_00000_11111_00000_00001_00000_11111_00000_11111_00000_00000_00010_11111_11111_11111_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b1010000101;  //node 645
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11111_00001_11111_00000_00000_00000_11111_00010_00001_11111_00010_11111_00000_11110_00000_00001_00000_11111_11111_11111_00001_00001_11111_11111_00000_11110_00000_11110_00000_00000_00010;

		#2
		WriteAddressSelect <= 10'b1010000110;  //node 646
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00000_00000_11111_00001_00000_00000_00001_11111_11111_00001_00001_11110_00001_11111_00001_00000_11110_00000_00000_00000_00000_11110_00000_00000_00000_00000_11110_00010_00001;

		#2
		WriteAddressSelect <= 10'b1010000111;  //node 647
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_11110_00000_00000_11111_00001_00000_11111_00000_00001_11111_00001_11111_00000_00001_11111_00001_00000_11110_00001_00000_11111_11110_00001_00000_00000_00001_00000_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010001000;  //node 648
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00001_00001_11111_00001_11111_11111_00000_00001_00000_11110_00001_00000_00010_00000_00000_11111_00001_00001_00001_00000_00000_00001_11111_00001_11111_11110_00001_11110_00010;

		#2
		WriteAddressSelect <= 10'b1010001001;  //node 649
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_11111_00001_00000_11111_00001_11111_00000_00001_11111_00001_00000_00001_00001_00001_11111_00001_00010_11111_11111_00000_00000_00001_00000_00001_00001_11111_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b1010001010;  //node 650
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11110_11110_00000_00000_00000_00001_00010_11111_00000_00010_11111_00000_00000_00000_00001_00000_00001_11111_00010_00001_00000_11111_11111_11111_11111_00000_00001_00000_00010_11110_00010;

		#2
		WriteAddressSelect <= 10'b1010001011;  //node 651
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11100_11111_11111_00000_00000_00000_00000_00000_00001_00000_11111_00001_00010_00001_00000_00000_11111_00010_00010_00000_00001_00001_00000_00000_11111_00010_00001_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010001100;  //node 652
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_00000_00000_11111_11111_00000_00001_11111_11111_00000_00010_11111_00001_00001_11110_11111_00010_11110_00010_00000_11111_00001_00000_11100_00000_00010_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010001101;  //node 653
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00001_00000_11111_00000_11111_00001_00001_00001_11110_11111_00010_11111_00010_00000_11111_11110_00010_11111_00001_00000_00000_00010_00010_11111_11110_00001_00001_00010_11110;

		#2
		WriteAddressSelect <= 10'b1010001110;  //node 654
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_11111_11111_00000_00001_11110_00001_00000_00000_11110_11111_00010_11111_00000_00001_11110_00000_11101_11111_00010_00000_00000_00001_00010_11110_00000_00010_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b1010001111;  //node 655
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_11110_11110_11111_11111_00010_11111_00001_00000_00000_00000_11111_00010_11111_00000_00010_11111_00000_00000_11110_11111_11111_00010_11111_11111_00010_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1010010000;  //node 656
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_00001_00000_00000_00000_00010_11111_00000_00000_00001_00000_11110_00001_11111_11111_00000_11110_00000_11110_00001_00001_00001_00001_00000_00000_11111_00010_00010_11111;

		#2
		WriteAddressSelect <= 10'b1010010001;  //node 657
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00011_11111_11110_00001_00001_11110_11111_00011_11111_00000_11110_00000_11110_11111_11111_11111_00010_11110_11110_00000_00000_00001_00001_11111_00000_00000_00001_00000_00010_11111_11111;

		#2
		WriteAddressSelect <= 10'b1010010010;  //node 658
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_00000_00000_11111_11111_00010_00000_00001_00010_00010_00010_11111_11111_00000_00000_00001_11111_11110_11110_11111_11110_11111_00001_11111_11111_11111_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b1010010011;  //node 659
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00010_00010_00001_00000_11110_00010_00001_11111_11111_00001_11111_00000_00000_11111_00001_00001_00000_00000_00000_11111_11111_00000_00000_00000_00000_11110_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b1010010100;  //node 660
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_11110_11111_11111_00000_00010_00000_11111_11110_11110_11111_11111_00001_11110_00000_11111_00010_11111_00000_00010_00000_11110_11110_00000_00001_00000_00001_11110_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1010010101;  //node 661
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00000_11110_00000_00001_11111_11111_00000_00000_00000_11111_00010_11111_11111_00000_00000_11111_00000_11111_00000_00010_00000_00001_11111_11111_00000_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010010110;  //node 662
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_00001_00001_11111_11111_11111_00000_00000_00000_00000_11111_11111_00001_00001_00000_00000_00000_11110_00000_00000_00000_11110_00000_11111_00010_00000_11111_11111_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b1010010111;  //node 663
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11111_11111_11110_00001_00000_00000_00000_00001_00000_00000_00000_00010_00000_00001_00000_00010_11111_00001_00001_11110_11111_00000_11111_11110_00000_00000_00000_11111_11110_11111;

		#2
		WriteAddressSelect <= 10'b1010011000;  //node 664
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00001_00001_11111_00001_11110_00010_00001_00001_11111_00001_00000_00000_00000_00010_00000_00000_00000_00100_11111_11111_11110_00000_00001_00000_11111_00000_11110_00000_00001_00001;

		#2
		WriteAddressSelect <= 10'b1010011001;  //node 665
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00000_00001_00001_00000_00010_00001_00000_00001_00000_00000_00001_00001_00000_00001_00000_00000_11111_00000_00001_11111_11111_11111_00001_11111_11110_00001_11110_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010011010;  //node 666
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_11111_00001_11111_00000_11111_00000_00001_00000_00000_11111_00000_00010_00000_11111_11111_00000_00001_11110_00000_11111_00001_11110_00010_00001_11111_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b1010011011;  //node 667
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_11111_00000_00000_00001_00000_00001_11110_11110_11110_11111_00010_00000_00000_00001_00000_11110_00001_00001_11111_11111_00000_00001_11111_00000_11110_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010011100;  //node 668
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_11111_11111_00000_00001_00000_00001_00000_00001_00001_00001_00001_11111_00001_11111_11111_11111_00001_00001_00001_00001_11111_00001_11111_00010_00001_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010011101;  //node 669
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00010_00000_00000_11111_00000_00000_00000_00000_11111_00000_00001_00001_00001_11110_00000_00001_00000_00001_11110_00000_11111_00010_11110_11111_11110_00000_00000_11111_00010;

		#2
		WriteAddressSelect <= 10'b1010011110;  //node 670
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_11111_00000_00001_00001_00000_00000_00001_11111_00001_00000_00001_11111_11111_00000_00010_00000_00000_00000_11110_00001_00000_11111_00010_00000_00000_00000_00000_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b1010011111;  //node 671
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_11111_00000_00001_00000_11111_00001_00000_11111_00000_11111_11111_00010_00000_11111_11111_11111_00000_00001_11111_11111_00001_11111_11110_11110_00001_11110_11111_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1010100000;  //node 672
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11110_00000_00001_11111_00001_00001_00001_00001_00001_00000_00001_00000_00001_11111_00000_00001_00001_00001_00000_00000_00001_00010_00000_00001_00001_00000_00010_00000_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1010100001;  //node 673
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_11111_00000_00000_00001_11111_00001_00000_11110_11111_00000_00000_00000_00010_00001_00001_11111_00001_00000_00000_00001_00000_11111_00000_11111_00001_11110_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1010100010;  //node 674
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11111_11111_00001_00001_00000_00000_11110_11111_00010_00001_00000_00001_00000_11111_11110_11111_00000_00000_11110_00000_00000_00000_00001_00000_00001_00000_11111_11111_00001_11111;

		#2
		WriteAddressSelect <= 10'b1010100011;  //node 675
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11111_00000_00000_00000_11111_00001_11111_00001_00000_00010_11110_11111_00001_00001_00001_00000_00000_00000_00000_00001_00010_11111_00000_00000_11110_11110_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b1010100100;  //node 676
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00001_00010_00001_00001_00010_11111_11111_00001_11111_00000_00000_11111_00001_00001_00000_00010_00001_00001_11111_00000_11110_00000_00010_11111_00000_00000_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1010100101;  //node 677
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_00001_00010_00010_00001_11111_00000_00010_00000_11111_00000_00001_11111_00000_11111_00000_00001_00001_00001_00000_00001_00000_11111_11111_00001_00000_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010100110;  //node 678
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00001_00001_00001_11111_00001_11111_00000_00000_11111_00001_00010_00000_00000_00000_00000_11111_00000_11111_00001_11111_00001_00001_11110_00000_00001_00010_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1010100111;  //node 679
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00001_00010_00001_11110_11110_00001_00001_00000_00000_00001_00010_11111_11111_00001_11111_00000_00010_00000_11111_00001_00001_00000_00000_00001_00000_00001_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010101000;  //node 680
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_11101_00001_00000_00001_00001_11110_11111_00000_11111_11111_00000_00000_00001_00000_00001_00000_11110_00000_00001_11111_00000_00001_11111_00000_11110_00000_00001_00010_00000_11111_11111;

		#2
		WriteAddressSelect <= 10'b1010101001;  //node 681
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11110_00000_00000_11111_11110_11111_00000_00000_11111_11111_00001_00001_11111_00001_00001_11110_11110_00010_00001_00010_00001_00001_00001_11111_00001_11111_00000_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b1010101010;  //node 682
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00001_11111_11111_11111_11111_00000_11110_00001_11111_00000_00010_00000_00010_11111_11110_00000_00001_00000_00010_00000_00001_11111_11110_00000_00001_00010_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b1010101011;  //node 683
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00001_11111_00001_11111_00000_00000_00001_00001_11111_00000_00001_11110_00000_00001_11110_00001_11111_00000_11111_00000_00000_00000_11111_11101_11111_00001_00001_00000_00010;

		#2
		WriteAddressSelect <= 10'b1010101100;  //node 684
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_00001_11111_00010_00000_00001_00010_00010_00001_00000_11111_00001_00000_00001_00001_11111_00000_00000_11111_00000_11111_00001_00000_00001_11111_11110_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1010101101;  //node 685
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00001_00001_00001_11110_00000_00000_00010_11110_11111_00001_11111_00000_11110_00010_00000_11111_00001_00000_11110_00000_11111_00000_00000_00000_11111_00000_00000_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010101110;  //node 686
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00000_11111_00001_11111_00000_11111_00010_11101_11110_11110_00001_11111_00000_11110_00000_00000_11110_11111_00000_00000_00001_00000_00000_00001_00010_00000_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1010101111;  //node 687
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00001_11111_00010_11110_00000_11111_00001_00000_11111_00001_00010_00010_11111_00010_00001_11110_11110_00000_00001_00000_00000_00000_11111_00001_11110_11111_11111_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b1010110000;  //node 688
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11111_00001_00000_11111_11111_11111_00001_00010_11111_00000_00000_00000_00000_00000_11110_00010_00001_11111_00001_00001_00000_00000_00000_00001_00000_00000_00000_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b1010110001;  //node 689
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_11110_00001_11111_00010_00000_00010_00010_00000_11111_00000_00001_00000_00001_00010_11110_00001_00000_11111_11111_00000_00010_11111_00001_11111_00000_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010110010;  //node 690
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00001_11110_00000_11110_00000_11110_00001_00000_11111_11111_00001_00000_00001_11111_00001_11110_00000_00000_00010_00000_00001_00001_00010_00001_11111_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b1010110011;  //node 691
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_00000_11111_00001_00001_11110_00000_00000_00001_00000_00001_00000_00001_00010_00001_11111_00000_11111_11111_11110_00001_11111_11111_00000_11111_11111_11110_11111_00001;

		#2
		WriteAddressSelect <= 10'b1010110100;  //node 692
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00010_11110_00000_11111_11111_00000_11111_00001_00000_11111_00000_11111_00000_00001_00001_00001_00000_11110_11111_00000_11111_00001_11110_11111_11111_11111_11111_11111_00001_11110;

		#2
		WriteAddressSelect <= 10'b1010110101;  //node 693
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_11111_00000_00001_00001_00001_11111_00000_00001_00000_00010_11111_11110_00001_00000_11111_00001_11111_11111_00000_11111_11110_00001_00000_00010_11111_00010_11110_00001;

		#2
		WriteAddressSelect <= 10'b1010110110;  //node 694
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00010_00000_00000_00000_11110_00001_00000_00000_00000_11111_11111_00000_11110_11111_00000_00001_11111_00000_00010_11111_11110_00000_00001_00001_11110_00001_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010110111;  //node 695
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00010_00000_00000_00000_00010_00000_00001_00000_00001_00000_00000_00010_00001_11111_00000_00011_00001_00000_11111_11111_11111_00000_11111_11111_00000_00010_00001_00000_00001_00010;

		#2
		WriteAddressSelect <= 10'b1010111000;  //node 696
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00010_00001_11111_11111_00000_00010_00001_00010_11111_00010_00000_00001_00001_00001_11111_00000_00000_00001_00000_00000_00000_00000_00001_00001_11111_11111_11111_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1010111001;  //node 697
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_00000_00010_11110_11111_11111_00000_11111_00010_00001_00010_11111_00010_00001_11111_11110_11111_00000_00000_00010_00000_11111_11110_00000_11111_11111_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b1010111010;  //node 698
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_11111_00010_00001_00001_00001_11111_00000_00000_11111_11111_00001_00001_11111_11110_00000_00010_00001_11111_11111_00001_00001_00000_00000_00000_00000_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010111011;  //node 699
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_11110_11111_00000_11110_00000_11111_11111_11111_11111_00001_00000_11111_00000_11110_00000_11111_00000_11111_00001_00001_00010_00010_00000_11110_00001_00001_00000_00000_11111_11110;

		#2
		WriteAddressSelect <= 10'b1010111100;  //node 700
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00000_11110_00000_00001_00000_00000_00001_11111_00000_11111_00000_00001_00000_00001_11111_00001_00000_00000_11110_00000_11111_00000_00000_00001_00001_00001_00010_11110_00010;

		#2
		WriteAddressSelect <= 10'b1010111101;  //node 701
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00001_00010_00010_11111_11111_00001_00000_11111_11110_00000_11110_11111_11111_00000_00000_11111_11111_00000_00000_00000_00000_11111_11111_00000_00010_11111_00000_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b1010111110;  //node 702
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_00001_00000_00001_00001_11111_00001_00000_00001_00001_00001_11110_00000_00000_11111_00000_00001_00001_11110_00001_11111_00001_00000_11111_11111_00000_00001_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1010111111;  //node 703
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11110_11111_00010_11111_00001_00001_00000_00010_00010_11111_11111_00000_00000_00001_00001_11111_00010_00000_00010_11111_00000_11111_00000_00000_00000_11111_11111_00000_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011000000;  //node 704
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_11110_00010_00000_00000_00001_11110_00010_00000_00000_00000_00000_00010_00001_11111_00001_00001_11111_11111_00000_00000_00001_00000_11111_00000_11111_11111_11111_00010_11110;

		#2
		WriteAddressSelect <= 10'b1011000001;  //node 705
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11111_11111_00001_00000_11111_11111_00000_00000_00001_11111_00000_11111_00001_11111_00010_00000_00000_00000_00001_00001_00010_00001_11111_11111_11111_00010_00000_11110_00000;

		#2
		WriteAddressSelect <= 10'b1011000010;  //node 706
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11110_00000_00000_00001_00001_00001_00001_11110_11110_00000_00001_00000_11111_00010_11111_00000_00001_00000_11110_00000_00010_00001_00000_00001_00000_00000_00001_00001_00000;

		#2
		WriteAddressSelect <= 10'b1011000011;  //node 707
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_00000_00000_00000_11111_11111_00001_11110_00000_00000_11111_00010_00001_11111_00000_11111_11111_00001_00000_00010_11111_11111_00001_11111_00000_00000_11111_11111_11111_00010;

		#2
		WriteAddressSelect <= 10'b1011000100;  //node 708
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_00000_00010_11111_00001_00000_11111_00000_00000_11110_00000_11111_00000_00000_00001_11111_11111_00010_00001_00000_11111_00000_11111_11111_00000_00000_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011000101;  //node 709
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_00001_00000_00000_00001_00000_00000_00000_00000_11111_00010_11111_00000_11111_00001_00000_00010_00000_00001_11111_00000_00000_11111_00001_00000_00001_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b1011000110;  //node 710
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_11111_11111_11110_11111_00001_11111_00000_11111_00000_00000_00001_00000_11111_00001_11111_00000_11111_00001_00000_00000_11111_00000_11111_11111_00000_00001_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011000111;  //node 711
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11110_00000_00000_00001_00001_11111_11110_00001_00000_00000_00001_00000_00000_11111_11110_00000_00001_00000_00001_00000_00001_00010_00001_11111_00000_00001_00000_11111_11111_11110;

		#2
		WriteAddressSelect <= 10'b1011001000;  //node 712
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00010_11111_00000_00000_00000_00001_00001_11111_00000_00000_00000_00000_11111_00001_00000_00001_11110_11111_00000_00001_00001_00000_00000_00000_00001_00000_11111_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b1011001001;  //node 713
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_11110_00000_00000_00000_11111_00000_11111_00001_11111_00001_00000_00000_11111_11111_11111_00000_00000_11111_11111_00000_00000_00001_00010_11111_00001_00000_11110_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011001010;  //node 714
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_00000_00000_11111_00000_00000_00000_11110_00001_00000_00001_11111_00000_00000_00010_11111_00000_11111_00010_00000_11111_00000_11110_11111_11111_00001_11111_11111_00001_11111_11111;

		#2
		WriteAddressSelect <= 10'b1011001011;  //node 715
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00010_11111_00000_00001_00000_00001_00000_00001_00000_00000_11111_00001_00010_00001_11111_00000_00001_00000_00001_00000_00001_00000_00000_00001_00000_11110_00001_00000_11110_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011001100;  //node 716
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00010_11111_00010_11111_00010_00000_00000_00000_11111_00001_11111_00000_00000_00000_00001_00001_00001_11111_00000_11110_00000_00000_00000_00001_11111_11111_00001_00001_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011001101;  //node 717
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00010_00000_00001_11110_00000_11111_00000_00000_11111_11111_00000_00000_00001_00010_00000_11111_00000_00001_11110_11111_11111_11111_00000_00010_11111_00001_00000_00000_11111_00001_00010;

		#2
		WriteAddressSelect <= 10'b1011001110;  //node 718
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_00000_00001_11111_00000_11111_00001_00001_00000_00000_11111_11111_00001_00001_11111_00010_11111_00000_11111_11111_00000_00000_11111_11111_00001_00001_00000_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b1011001111;  //node 719
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_11110_11111_11111_00000_00000_11111_00001_11111_00000_11111_00000_11111_00000_11111_11111_00001_11110_00000_00001_11110_11111_00000_00010_11111_00000_00000_00001_00001_00001;

		#2
		WriteAddressSelect <= 10'b1011010000;  //node 720
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00010_00001_00000_00001_11111_00000_00001_11110_00000_11111_00000_00010_00000_00000_00000_00001_00000_00000_00000_11111_11111_11110_00000_11110_00001_00000_11110_11111_11111_11111;

		#2
		WriteAddressSelect <= 10'b1011010001;  //node 721
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00001_00001_00000_00000_00001_00000_11110_00000_11111_00001_00000_11111_00010_11111_00001_11111_11111_11110_00001_11111_11111_00001_00000_00000_00000_00001_00000_00001_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011010010;  //node 722
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00010_00001_11111_00000_00000_00000_00001_00000_00001_11111_00000_00001_00000_00001_11110_00000_00001_00000_00001_00001_00001_00000_11111_11111_00000_00000_00001_11111_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011010011;  //node 723
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_00000_11111_11111_11111_00001_00000_11111_11111_11111_00000_00000_11110_11111_00000_00000_11110_00000_11111_00000_00000_00000_00000_00001_00000_00000_00001_11111_00000_00010;

		#2
		WriteAddressSelect <= 10'b1011010100;  //node 724
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_11111_00000_00000_00001_00000_00010_00001_00000_11111_00000_00001_11111_00000_11111_11111_00001_00000_00000_00001_00001_11111_00010_00000_00001_00001_00001_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011010101;  //node 725
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00000_11110_11111_00000_11111_00010_11110_00000_00000_11111_00010_00001_00000_00000_00000_00000_00000_00010_11111_00000_00000_11110_00000_00001_00001_11110_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b1011010110;  //node 726
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_00010_00001_00000_00000_00000_00000_00001_00001_00000_00000_00000_00000_11111_00000_00001_00000_00001_00001_00010_11110_00000_00000_00001_11111_00001_11110_00000_11110_11111;

		#2
		WriteAddressSelect <= 10'b1011010111;  //node 727
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00000_00001_11111_00000_00001_00010_00001_11110_00000_00000_00000_00010_00010_00001_11110_11110_00000_11110_00000_11111_11110_00000_00001_00001_00001_11111_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011011000;  //node 728
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_11110_00000_00010_00001_11110_11111_00001_11111_11111_00001_00000_00000_00000_00000_00000_00010_11111_11111_11111_00000_00000_11111_00001_11111_11111_00000_00000_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011011001;  //node 729
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_11111_00000_00000_00001_11111_00000_00001_00000_00001_00010_00001_00000_00000_00000_00001_00000_00001_00001_11111_11111_11111_00000_00000_00001_00000_00001_11110_00001_11111;

		#2
		WriteAddressSelect <= 10'b1011011010;  //node 730
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_11111_00000_00001_00010_11111_00000_11111_11111_11111_00001_11111_00000_11111_00001_00001_00001_00000_00000_11111_00001_00000_00001_00000_00001_11111_11111_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011011011;  //node 731
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_11111_00000_00000_00000_11111_00000_11111_11111_11111_00000_11111_00000_00000_00000_00010_11111_11111_00001_00010_00000_00000_00001_11111_00000_00001_00001_11111_00001_00001_00010;

		#2
		WriteAddressSelect <= 10'b1011011100;  //node 732
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_00001_00000_00000_00001_00001_00000_00000_11111_00000_00000_11111_00000_11111_11111_11111_11111_11110_00001_00000_00001_11110_00010_00000_00001_11111_11110_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011011101;  //node 733
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00010_00010_00000_00001_00010_11111_11111_00001_00001_00001_00000_00001_11111_00000_00001_00001_00000_00001_00010_00000_00001_00001_11111_00000_00001_11111_00001_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b1011011110;  //node 734
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00001_00000_00000_00000_00000_00001_00001_00001_00001_00000_11111_11110_00001_00000_00000_00010_00001_00000_11111_11111_00001_11111_00000_11110_00000_00000_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011011111;  //node 735
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_11110_00000_11111_00001_11111_00000_00000_00001_00001_00010_00001_11111_11111_00001_00000_11111_00000_00001_00001_00000_00000_00000_00000_00000_00000_11111_00000_11111_00010;

		#2
		WriteAddressSelect <= 10'b1011100000;  //node 736
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11110_11111_00000_11111_00001_11111_00010_11111_00001_11111_00001_00001_00000_00001_11111_00001_00001_00000_00000_11110_11111_11111_11111_11111_00001_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011100001;  //node 737
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_11111_00010_00000_00000_00001_00000_00010_11111_11111_00001_00000_00000_11111_11110_00001_11111_00000_11111_00001_00000_00000_00000_11110_00010_11110_00001_11110_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011100010;  //node 738
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00010_00000_11111_00000_11111_00000_00000_00001_00000_00000_11111_00000_00000_00000_11111_00010_00000_00000_00001_11111_00000_11111_00001_00000_00010_11111_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011100011;  //node 739
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00000_00010_00000_11110_00010_00000_00000_00000_00001_00001_00000_00000_00000_00001_11110_00010_00001_00000_11111_00001_00001_00001_11111_11110_11111_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011100100;  //node 740
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00000_00000_00000_00000_11111_00000_00000_00001_11110_00001_00001_00001_00001_00000_00000_11110_00000_11111_00000_00000_11111_00000_00001_00000_11111_00000_00000_00001_00000_11110;

		#2
		WriteAddressSelect <= 10'b1011100101;  //node 741
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00001_00001_00001_00000_11111_00001_11111_00000_11111_00000_00010_00000_00000_11110_00001_00000_00000_00000_11111_00010_11111_00001_00001_00000_11111_00001_11111_11111_00010_00000;

		#2
		WriteAddressSelect <= 10'b1011100110;  //node 742
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_11111_00010_11111_00000_00000_00001_11111_00000_00000_00000_11111_00001_00000_00000_00000_00001_00010_00000_00000_00000_00000_11111_00001_11111_00000_11110_11110_11111_11110_00000;

		#2
		WriteAddressSelect <= 10'b1011100111;  //node 743
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00000_00010_11111_00001_00001_11111_00000_00000_00001_11110_11110_11111_11111_00000_00010_00000_11111_00010_00000_00001_00001_11111_00000_11111_00001_00000_00010_00000_00010_00000;

		#2
		WriteAddressSelect <= 10'b1011101000;  //node 744
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_11111_00000_00000_00001_11111_11111_11110_11111_11110_11111_00001_00000_00000_00000_00010_00000_11111_00000_00010_00000_00001_00001_11111_00000_11111_00001_00010_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011101001;  //node 745
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00001_11111_11111_11111_00000_00000_00000_11110_11111_00000_11111_00001_11111_11111_00001_11111_11110_11111_11111_00000_00000_00010_11111_00000_00001_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011101010;  //node 746
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_11111_00000_00000_00000_00000_11110_00010_00000_00000_11111_11111_00001_00000_00000_00000_00000_00001_00001_00001_00001_11111_00000_00000_00010_00001_11111_11111_00000_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011101011;  //node 747
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00001_11110_00001_00000_11111_00010_00001_00000_11110_00000_00001_11111_00000_11111_11111_00000_00000_11111_00001_11111_11111_11111_00000_00000_11111_00000_00000_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011101100;  //node 748
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00000_00001_11111_00000_00010_00001_11111_11111_00000_11111_00000_11111_00001_11111_00001_00001_11111_00001_00000_00000_00001_11110_11111_11111_00000_00010_00000_00001_00001_11111;

		#2
		WriteAddressSelect <= 10'b1011101101;  //node 749
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_11111_11111_11110_00000_00000_11110_00010_00010_00000_00000_11111_11111_00001_00010_11111_11111_00000_00000_00000_00000_00010_00000_00000_00001_00000_00010_11111_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011101110;  //node 750
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00000_00010_00001_00000_00001_00000_00010_00000_11111_00001_00000_11111_11111_00000_00001_11111_00000_11111_11111_11111_00000_00000_00000_00001_00001_11111_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1011101111;  //node 751
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11110_00000_11111_00001_00001_11111_00001_00000_00001_11110_11111_00001_11110_11111_00001_00000_11111_11111_00000_11111_00000_00000_00000_00010_00001_00001_00000_00001_00000_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011110000;  //node 752
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00000_11111_00001_00000_00001_00001_00000_00000_11111_00000_00000_00000_00001_00001_00001_00001_00000_00001_11111_00000_00000_00000_00001_00000_00000_11110_00001_00001_00010_00000;

		#2
		WriteAddressSelect <= 10'b1011110001;  //node 753
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_00010_00000_11110_00000_00000_00001_00000_11111_11111_00000_00001_11111_00000_11111_00000_00000_00001_00000_00001_00010_00001_00000_00000_00001_00001_00010_00001_00000;

		#2
		WriteAddressSelect <= 10'b1011110010;  //node 754
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00000_00000_00000_11111_00000_00000_00010_00000_11111_00001_11110_00010_11111_00000_11110_11111_00001_11111_11110_11110_00000_00000_00010_00000_00000_00001_00000_00001_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011110011;  //node 755
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11110_11110_11111_00001_11111_00010_00001_00001_00000_11111_00000_00001_00000_11110_00001_00000_00000_00001_00001_00000_00001_00000_00000_00010_11110_00001_00010_00000_00000_00010;

		#2
		WriteAddressSelect <= 10'b1011110100;  //node 756
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00001_11111_00001_00000_00001_00000_11110_11110_00001_00000_00001_00000_00000_11111_00001_00000_11110_00000_11111_00001_00000_11110_00010_00000_11111_00001_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011110101;  //node 757
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00000_00001_00010_11111_00000_11111_00010_11111_11110_00000_00000_00000_11111_11111_00010_00001_00001_11111_00000_00000_00000_00000_11111_11110_00001_00000_11111_11111_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011110110;  //node 758
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00001_11111_00000_11111_00000_00000_11111_00000_11111_00000_00001_00000_00010_00000_00000_00010_00001_00010_11111_00001_11110_00001_00001_00000_00000_11111_00001_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1011110111;  //node 759
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00000_00000_00001_00000_11111_00000_00000_11111_00000_00001_00000_11111_00000_00000_00001_00000_11111_11110_00001_00000_00001_00001_00000_00001_00000_11111_00000_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011111000;  //node 760
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00001_00000_00000_00010_11110_11111_00001_11111_11111_11111_00000_00000_11111_11111_11111_00001_00000_00001_00000_11111_11111_00000_00000_00001_00010_00000_00000_00001_00001_11111_00001;

		#2
		WriteAddressSelect <= 10'b1011111001;  //node 761
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_11111_00000_11111_11111_00000_00000_11110_11110_00001_00000_11111_00000_00000_00000_00000_00001_00000_00001_11111_00001_11111_11111_11111_00001_11111_11111_00001_00001_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011111010;  //node 762
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_11111_00000_00000_11111_00001_00000_00000_00010_00000_00000_00000_00000_11110_00010_11111_00010_00010_00001_00000_11111_00000_11110_11111_00010_11111_00001_11111_00000_00000;

		#2
		WriteAddressSelect <= 10'b1011111011;  //node 763
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00000_00000_00000_11111_11111_00001_00010_11110_00000_00000_00000_00000_00001_00001_00000_00001_11111_00001_00001_00000_11110_00001_11111_00010_00000_00001_00010_00001_00001;

		#2
		WriteAddressSelect <= 10'b1011111100;  //node 764
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00001_00010_00000_00000_00001_00000_11110_00000_00000_11110_11110_00000_00001_00001_11111_00000_11110_00010_11111_11111_00000_00010_00001_00001_00001_00001_00001_00010_11111_00001_00001;

		#2
		WriteAddressSelect <= 10'b1011111101;  //node 765
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_11111_11111_11111_11111_00000_00000_00000_11110_00000_00000_00000_11111_00001_00010_00000_11111_00000_00000_00000_00001_00001_00010_11111_00000_00001_11110_00000_00000_00000_00010;

		#2
		WriteAddressSelect <= 10'b1011111110;  //node 766
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00001_11111_11110_11110_00000_00000_11111_00001_00001_00000_00000_11111_00000_11111_00000_11111_00000_00000_00000_00000_11111_00001_00000_00000_11110_11111_00001_00000_00001;

		#2
		WriteAddressSelect <= 10'b1011111111;  //node 767
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_11111_00000_11111_00000_00000_00000_11111_00001_00001_11110_00000_00000_00001_00001_00001_00010_00000_11111_11111_00001_11111_11111_11111_00010_00000_11111_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1100000000;  //node 768
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00001_00000_00000_11110_00001_00000_00000_00000_00001_00000_00001_00001_00000_11111_00010_00001_00001_00000_00001_00000_00001_00000_00001_00000_11111_00001_11111_00001_11111_11111_00001;

		#2
		WriteAddressSelect <= 10'b1100000001;  //node 769
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00010_00001_00010_00001_00001_00000_11110_00000_11111_11111_00000_00000_00001_00010_00010_00000_00000_00000_00000_00001_00001_00010_11111_00000_00001_11111_00001_00010_00001_11110_11111_11110;

		#2
		WriteAddressSelect <= 10'b1100000010;  //node 770
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_00010_00001_00000_00000_00001_00000_11111_11111_00010_00001_11111_00000_00001_00000_11111_11110_00000_00001_11111_00001_00001_00000_00000_11110_00000_00001_00000_00010_11111_00001;

		#2
		WriteAddressSelect <= 10'b1100000011;  //node 771
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_11111_11111_00001_00001_11110_11111_00001_11110_11111_00000_11111_00000_00010_00000_00000_00000_00000_00000_11110_11111_11111_00001_00000_00001_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1100000100;  //node 772
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_11111_11111_00000_11111_00000_00001_00001_11111_00001_00000_11111_11111_11111_11111_00000_11111_11111_00000_11111_00000_00000_00001_00001_00000_00000_00000_00000_00001_11111_00000;

		#2
		WriteAddressSelect <= 10'b1100000101;  //node 773
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_00000_11111_00001_11111_00000_00001_11111_00001_00001_00000_00010_00000_11111_00010_00010_00001_00001_00000_00001_00001_11111_11111_11111_11111_00001_00000_11111_00000_00001_11110;

		#2
		WriteAddressSelect <= 10'b1100000110;  //node 774
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_00000_00001_00001_00010_00000_00000_00010_00000_00000_00001_00000_00001_00001_00001_00000_11111_00001_00001_00010_00000_11111_11111_11111_00000_00001_00010_00000_00000_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1100000111;  //node 775
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_00010_00000_11110_00010_00000_00000_11111_11111_00000_00000_11111_00000_00001_11110_00001_00001_00000_00001_00001_11111_11111_00010_11111_00000_00000_00010_00000_00000_00000_11110;

		#2
		WriteAddressSelect <= 10'b1100001000;  //node 776
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11111_11110_00000_00000_00001_11111_11111_11110_11111_11111_00001_00001_00001_00001_11111_00000_11111_11111_00001_11111_11111_00000_11111_00000_00000_00000_00001_11111_00000_11111_00000;

		#2
		WriteAddressSelect <= 10'b1100001001;  //node 777
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11111_11110_00000_00000_00000_11111_11111_11110_00001_11111_00010_00001_00001_11111_00010_00010_11111_00000_00000_00000_00010_00001_00000_00000_00001_00000_00000_00000_00000_00000_00000_11111;

		#2
		WriteAddressSelect <= 10'b1100001010;  //node 778
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_11111_00001_00000_00000_00000_00001_00010_11110_00000_11110_11111_00000_00000_00000_11111_11110_00000_00000_00000_11111_00010_00000_11110_00000_00000_11111_00000_11111_00000_00001_11111;

		#2
		WriteAddressSelect <= 10'b1100001011;  //node 779
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00001_00010_11111_11111_00000_00000_00001_11111_00001_00000_11110_00000_11111_00000_00001_00000_00000_00000_00000_11111_00000_00001_00000_00000_00001_00000_11111_11110_11110_00000_00001;

		#2
		WriteAddressSelect <= 10'b1100001100;  //node 780
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_11111_11111_00001_00001_00001_11111_00000_00000_00001_00000_00001_11111_11111_00001_00010_00001_00001_00000_00000_11110_11111_00010_11111_00000_00001_11111_00010_00010_11110_11111_11111;

		#2
		WriteAddressSelect <= 10'b1100001101;  //node 781
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b11110_00000_00010_00001_11111_11111_00000_00000_00001_00000_00001_00000_11111_00001_11111_00001_00000_00000_11111_11111_00010_11110_00001_11111_11111_00000_00001_00000_00000_00001_11110_00000;

		#2
		WriteAddressSelect <= 10'b1100001110;  //node 782
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00001_00000_00001_00000_00010_11111_00000_11111_11111_00000_00000_00000_11111_11111_11111_00000_00010_00000_11111_00000_11111_11110_00001_00000_00000_00000_00000_00001_11111_00000_00001_00000;

		#2
		WriteAddressSelect <= 10'b1100001111;  //node 783
		weightWriteEnable <= 1;
		#1
		writeIn <= 160'b00000_00000_11111_00000_00000_00001_00001_00000_11111_00000_11111_00000_11111_11111_11111_00001_00000_11110_00000_00001_11110_00000_11111_00000_00001_00000_11111_00000_00001_11110_11111_00001;


		#1
		weightWriteEnable <= 0;

		//Layer 1 Biases
		#2
		biasWriteEnable <= 1;
		#1;
		writeIn <= 160'b00000_00101_00000_00000_00010_11110_00100_00001_00000_00010_11111_00010_00000_11110_11110_11110_00010_11111_11100_00010_00000_00010_00001_10101_00010_00000_10110_11111_00010_00000_11110_00000;
		#1
		biasWriteEnable <= 0;



		//Layer 2 Weights
		#1
		LayerWriteSelect = 1;
		#1
		#2
		WriteAddressSelect <= 10'b0;  //node 0
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000101_111110_101101_111110_000011_000101_000010_000001_111111_000110;

		#2
		WriteAddressSelect <= 10'b1;  //node 1
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000100_000001_001110_000010_111000_000001_001101_111011_111101_110110;

		#2
		WriteAddressSelect <= 10'b10;  //node 2
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000010_111100_111110_000100_111110_111110_111010_000111_000110_000011;

		#2
		WriteAddressSelect <= 10'b11;  //node 3
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111110_001010_000010_110001_000101_111000_000111_000101_000000_000010;

		#2
		WriteAddressSelect <= 10'b100;  //node 4
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000000_111101_000000_110110_001010_111111_111110_001000_111000_111111;

		#2
		WriteAddressSelect <= 10'b101;  //node 5
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111110_000101_000101_000001_000011_101110_111100_000011_111111_000101;

		#2
		WriteAddressSelect <= 10'b110;  //node 6
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111010_000100_111011_001010_000010_111110_111010_111110_000110_111111;

		#2
		WriteAddressSelect <= 10'b111;  //node 7
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111100_000000_001100_111110_000111_000011_111010_111010_110111_000011;

		#2
		WriteAddressSelect <= 10'b1000;  //node 8
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b001010_110111_111000_111101_000000_000010_001010_111110_000101_000010;

		#2
		WriteAddressSelect <= 10'b1001;  //node 9
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000110_000001_000000_000111_111100_001001_111110_111100_110010_000110;

		#2
		WriteAddressSelect <= 10'b1010;  //node 10
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b110111_111100_111001_001000_000011_001000_111100_111011_000011_001101;

		#2
		WriteAddressSelect <= 10'b1011;  //node 11
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111000_111110_000111_000011_111100_111110_111100_001110_111010_000111;

		#2
		WriteAddressSelect <= 10'b1100;  //node 12
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111111_001001_000101_110100_001010_111110_111010_000010_111100_000110;

		#2
		WriteAddressSelect <= 10'b1101;  //node 13
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000010_000000_001001_000010_111111_000011_111000_000010_000011_110010;

		#2
		WriteAddressSelect <= 10'b1110;  //node 14
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b110110_111111_111111_000110_000011_000100_111001_110111_001000_001010;

		#2
		WriteAddressSelect <= 10'b1111;  //node 15
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b001000_111110_001010_000010_101000_000011_000101_111111_000110_111110;

		#2
		WriteAddressSelect <= 10'b10000;  //node 16
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111111_000111_111111_110101_001110_000100_000010_000001_111110_110110;

		#2
		WriteAddressSelect <= 10'b10001;  //node 17
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111010_001000_001110_001011_111001_111011_111110_010100_110111_110011;

		#2
		WriteAddressSelect <= 10'b10010;  //node 18
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111110_110100_111110_111010_110100_010000_001011_111110_000101_000011;

		#2
		WriteAddressSelect <= 10'b10011;  //node 19
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111001_000010_111110_000010_000010_001010_000111_111000_000100_110101;

		#2
		WriteAddressSelect <= 10'b10100;  //node 20
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111011_111001_111110_000010_110011_001110_000011_000101_000010_000110;

		#2
		WriteAddressSelect <= 10'b10101;  //node 21
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111111_111110_000001_111100_111000_001011_111000_000100_111110_000101;

		#2
		WriteAddressSelect <= 10'b10110;  //node 22
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000010_111110_111010_001010_000001_111101_000101_000110_111111_111110;

		#2
		WriteAddressSelect <= 10'b10111;  //node 23
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111100_000011_111101_000101_001000_000010_111101_000000_110000_001011;

		#2
		WriteAddressSelect <= 10'b11000;  //node 24
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111101_111101_000110_111100_001011_111010_111110_111010_001000_111100;

		#2
		WriteAddressSelect <= 10'b11001;  //node 25
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000011_000110_000100_000000_000001_110010_111010_000110_111010_000000;

		#2
		WriteAddressSelect <= 10'b11010;  //node 26
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000110_000101_111111_000100_000011_111010_000111_000110_101111_111001;

		#2
		WriteAddressSelect <= 10'b11011;  //node 27
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111110_010011_111101_111101_111110_000010_000010_111111_111101_111100;

		#2
		WriteAddressSelect <= 10'b11100;  //node 28
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000101_111111_111000_000110_110011_001101_000001_111011_111110_111101;

		#2
		WriteAddressSelect <= 10'b11101;  //node 29
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b111011_000010_111111_111000_111110_000010_000111_000101_000111_111010;

		#2
		WriteAddressSelect <= 10'b11110;  //node 30
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000100_111101_000001_000010_111010_000010_110101_111110_000111_001010;

		#2
		WriteAddressSelect <= 10'b11111;  //node 31
		weightWriteEnable <= 1;
		#1
		writeIn <= 60'b000000_111111_000001_111110_111110_111111_111110_000110_111110_000110;


		#1
		weightWriteEnable <= 0;

		//Layer 2 Biases
		#2
		biasWriteEnable <= 1;
		#1;
		writeIn <= 60'b00000_00101_00000_00000_00010_11110_00100_00001_00000_00010_11111_00010_00000_11110_11110_11110_00010_11111_11100_00010_00000_00010_00001_10101_00010_00000_10110_11111_00010_00000_11110_00000;
		#1
		biasWriteEnable <= 0;

		//=================================
		//--Reset Network--
		//=================================
		
		#2
		reset <= 1;
		#2
		reset <= 0;

		//=================================
		//--Define Input Vectors--
		//=================================

		//Input 0
		inputVectors[0] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000001100000000000000000000000000110000000000000111100000000011000000000000111110000000001100000000001111110000000000110000000001110000000000000011000000001110000000000000001100000111110000000000000000110001111100000000000000000011001111000000000000000000001111110000000000000000000000111100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 1
		inputVectors[1] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000111110000000000111100000000111111000000000011100000001111111100000000001100000011111100110000000001110000011111100011000000000111000011111000001110000000011100111110000000111000000001111111110000000011100000000011111100000000001110000000000010000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000;
		//Input 2
		inputVectors[2] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000001111110000000000000000000111111100000000000000000011111110000000000000000001111110000000000000000000111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 3
		inputVectors[3] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000111111111110000000000000001111111111111100000000000001111110000001110000000000001111110000000111100000000001111110000000111110000000011111111000000011111000000001111111000000001111000000000111111000000001111100000000000011100000001111100000000000000111000000111110000000000000011110000111110000000000000000111111111111000000000000000000111111110000000000000000000001111100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 4
		inputVectors[4] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111100000000000000000001110000110000000000000000011100000001000000000000000111100000000100000000000000000000000000010000000000000000000000000001000000000000000000000000001100000000000000000000000000110000000000000000000000000011101011100000000000000001111111111100000000000000011111111111100000000000100111111000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 5
		inputVectors[5] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000011111111000000000000000001111111111000000000000001111111111000000000000000011111111100000000000000000111111110000000000000000000111111000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 6
		inputVectors[6] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000001111111000000000000000000001110001110000000000000000001110000111000000000000000000110000001100000000000000000000000000110000000000000000000000000011000000111000000000000000001100011111110000000000000001100111111111000000000000000111111100001000000000000000111110000001100000000000000011110000000100000000000000111100000000000000000000001111000000000000000000000001110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 7
		inputVectors[7] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001111111000000000000000000001111011110000000000000000001111000011100000000000000001111100001110000000000000000111110001110000000000000000000111111110000000000000000000001111110000000000000000000000011111110000000000000000000000111111100000000000000000000000001111100000000000000000000000001111000000000000000000000000000111000000000000000000000000001111000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 8
		inputVectors[8] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111100000000000000000000011111111000000000000000000011100011100000000000000000011100001110000000000000000000000000111000000000000000000000000001110000000000000000000000000111111000000000000111000000011111110000000000011100000001111111000000000001110000000111011110000000001111000000011111110000000000111000000001111111000000000011100000000111111000000000001110000000000111000000000000111000000000000000000000000011100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 9
		inputVectors[9] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111100000000000000000000000111111000000001100000000000111001100000011111000000000011101110000111111000000000011100111000111111000000000001110011100111110000000000000110001111111110000000000000111000111111100000000000000011100011111100000000000000001111101111000000000000000000011001111000000000000000000001110111100000000000000000000111111100000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 10
		inputVectors[10] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000001111111111111000000000001111111000000001110000000001111100000000000111000000000111000000000000011100000000011000000000000001110000000001100000000000000111000000000110000000000000011100000000111000000000000001110000000001100000000000001110000000000110000000000000111000000000011100000000000111000000000001111000000000111100000000000011111000001111000000000000000111111111111000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 11
		inputVectors[11] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000011111111111100000000000001111111000000111000000000011111100000000001100000000011100000000011000011000000001100000000111110001100000000100000000111111100110000000000000000011100010111000000000000000011100001011100000000000000011100000001100000000000000001110000001110000000000000000110000000110000000000000000011000000110000000000000000001100000110000000000000000000111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 12
		inputVectors[12] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111100000000000000000000011111110000000000000000000011100011000000000000000000011100001100000000000000000011100000110000000110000000001100000011000111111100000000110000011011111110000000000011000011111111000000000000001100011111110000000000000000010111111000000000000000000001111100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 13
		inputVectors[13] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111000000000000000001111111111111000000000000001111110000011110000000000001111100000000001100000000001111000000000000110000000000111000000000000001100000000111000000000000000010000000011100000000000000011000000001111000000000000001100000000111100000000000001100000000011111100000000011110000000000111111000000111110000000000000011111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 14
		inputVectors[14] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111111111111111111000000001111111111111111111000000000111111111111111111000000000000100111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 15
		inputVectors[15] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000011000000000011110011100000001110000000001111111100000000011000000000110000110000000001100000000011000010000000000110000000011000001000000000011000000001100000110000000001100000000110000011000000000110000000011000000100000000011000000001000000011000000001000000000100000000100000000100000000010000000011000000110000000000000000000110000011000000000000000000001100011000000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 16
		inputVectors[16] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111111000000000000000000011110000110000000000000000011100000011000000000000000001100000000100000000000000001100000000110000000000000000110000000011000000000000000011000000001100000011000000001100000000100011111100000000011000000111111111110000000000100001111111110000000000000000111111110000000000000000000111111000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 17
		inputVectors[17] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000011100000000111000000000000011110000000001100000000000111110000000000110000000000111110000000000011000000001111100000000000001110000001111100000000000000011000001111000000000000000001110011111000000000000000000111111110000000000000000000011111110000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 18
		inputVectors[18] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111100000000000000000000011111111000000000000000000001111000000000000000000000001111000000000000000000000000111000001100011000000000000001100001111001111000000000000111000011100011110000000000001110001110000011000000000000011100111000001110000000000001111111100000011000000000000011111110000001100000000000000111111000000111000000000000000011100000011000000000000000000111000001100000000000000000011100000110000000000000000000111000111000000000000000000011110011100000000000000000000111111100000000000000000000001111110000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		//Input 19
		inputVectors[19] <= 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000111111100000000000000000001111000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000110000000000000000001111111111100000000000001111111110000000000000011111111001100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
