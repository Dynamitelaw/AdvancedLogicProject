/*
 * This file describes the behaviour and IO of Layer 1. 
 * All modules needed for Layer 1 are instantiated here.
 */

`include "GlobalVariables.v"


module Layer1_Controller (
	//Inputs
		reset,
		//Timing
		clk, inputsReady, queueEmpty, outputsRecieved,
		//Memory updating
		weightWriteEnable, biasWriteEnable, WriteAddressSelect, writeIn, 
		//Data
		queueOut,

	//Outputs
		//Timing
		outputsReady, dequeue,
		//Data
		layer1Output
	);

	//Inputs
	input reset;
	input clk;
	input inputsReady;
	input queueEmpty;
	input outputsRecieved;

	input weightWriteEnable;
	input biasWriteEnable;
	input [9:0] WriteAddressSelect;
	input [`RELU_NODES*`LAYER_1_BIT_WIDTH-1:0] writeIn; 

	input [9:0] queueOut;

	//Outputs
	output outputsReady;
	reg outputsReady = `FALSE;

	output dequeue;
	reg dequeue = 0;

	output [`RELU_NODES*`LAYER_2_IN_BIT_WIDTH-1:0] layer1Output;
	reg [`RELU_NODES*`LAYER_2_IN_BIT_WIDTH-1:0] layer1Output;  //buffer layer1Output to allow for async pipeline

	//Internal variables
	reg processFinished = `FALSE;
	reg idle = `TRUE;


	//--Instantiate modules--

	reg [9:0] nodeAddress;
	wire [`RELU_NODES*`LAYER_1_BIT_WIDTH-1:0] weightStorageBus;
	Layer1WeightStorage weightStorage(
		//Inputs
		.writeEnable(weightWriteEnable), .NodeSelect(nodeAddress), .writeIn(writeIn), 
		//Outputs
		.readOut(weightStorageBus)
	);

	reg wBuffer_A_Write = `FALSE;
	wire [`RELU_NODES*`LAYER_1_BIT_WIDTH-1:0] wBuffer_A_Out;
	NodeWeightBank weightBuffer_A(
		//Inputs
		.writeEnable(wBuffer_A_Write), .writeIn(weightStorageBus), 
		//Outputs
		.readOut(wBuffer_A_Out)
	);

	reg pstoreReset = `TRUE;
	wire [`RELU_NODES*`LAYER_1_OUT_BIT_WIDTH-1:0] pstoreOutput;
	pStore plusStore(
		//Inputs
		.clk(clk), .clr(pstoreReset), .weightsIn(wBuffer_A_Out), .biasesIn(writeIn), .biasWriteEnable(biasWriteEnable),
		//Outputs
		.sumOut(pstoreOutput)
	);

	reg reluTrigger = `FALSE;
	wire [`RELU_NODES*`LAYER_2_IN_BIT_WIDTH-1:0] reluOutput;
	RELU relu(
		//Inputs
		.sumIn(pstoreOutput), .trigger(reluTrigger),
		//Outputs
		.layer1Out(reluOutput)
	);


	//--Controller behaviour--

	always @(posedge clk or posedge reset or posedge queueEmpty or posedge idle) begin : Layer1_proc
		//---------------------------------------
		// Async reset
		//---------------------------------------
		if (reset) begin
			outputsReady <= `FALSE;
			processFinished <= `FALSE;
			idle <= `TRUE;
			wBuffer_A_Write <= `FALSE;
			pstoreReset <= `TRUE;
			reluTrigger <= `FALSE;
		end

		//---------------------------------------
		// Idle processing and wakeup
		//---------------------------------------

		else if (idle) begin
			//Wake up from idle if we have something we can process
			if ((inputsReady == `TRUE) && (queueEmpty == `FALSE) && (outputsReady == `FALSE)) begin
				//The input layer is ready, and the output buffer of layer1 is empty. Ready to process
				processFinished <= `FALSE;
				idle <= `FALSE;
				wBuffer_A_Write <= `TRUE;
				pstoreReset <= `FALSE;  //enable pstore
				//reluTrigger <= `FALSE;
			end

			if ((outputsReady == `TRUE) && (outputsRecieved == `TRUE)) begin
				//The next stage has recieved our outputs
				outputsReady <= `FALSE;
			end
		end

		//---------------------------------------
		// Steady-state and near-end processes
		//---------------------------------------

		else begin
			//The input queue is empty. Near end of processing stage
			if (queueEmpty) begin
				//Turn off buffer writes. 
				wBuffer_A_Write <= `FALSE;
				// wBuffer_B_Write <= `FALSE;

				if (processFinished == `TRUE) begin
					//The input image has been processed by this stage

					layer1Output <= reluOutput;  //Store output of RELU to output buffer
					reluTrigger <= `FALSE;  

					outputsReady <= `TRUE;  //Notify next pipeline stage
					pstoreReset <= `TRUE;  //reset pstore

					idle <= `TRUE;  //go into idle state
				end
			end

			//Steady-state Positive clock edge events
			if ((queueEmpty == `TRUE) && (processFinished == `FALSE)) begin
				//This is the last pixel to be added. Get ready to shut down this pipeline stage
				reluTrigger <= `TRUE;
				processFinished <= `TRUE;
			end
		end
	end
	

	//---------------------------------------
	// Constant processes
	//---------------------------------------

	//Dequeue control
	always @(inputsReady or queueEmpty or clk) begin : dequeue_proc
		dequeue = inputsReady && (~queueEmpty) && clk && (~outputsReady);
	end
		
	//MUX for weightStorage address
	always @(weightWriteEnable or biasWriteEnable or queueOut or WriteAddressSelect) begin : address_mux
		if ((weightWriteEnable) || (biasWriteEnable)) begin
			nodeAddress <= WriteAddressSelect;
		end
		else begin
			nodeAddress <= queueOut;
		end
	end

endmodule
