
module multStore ( clk, clr, layer2In, weightsIn, biasesIn, biasWriteEnable, 
        sumOut );
  input [3:0] layer2In;
  input [59:0] weightsIn;
  input [59:0] biasesIn;
  output [99:0] sumOut;
  input clk, clr, biasWriteEnable;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n192, n193, n194, n195, n196, n198,
         n199, n200, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n225, n226, n227, n228, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n280,
         n281, n282, n283, n284, n285, n286, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n410, n411, n412, n413, n414, n415, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n430, n431, n432, n433,
         n434, n435, n436, n437, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n842, n843, n844, n845, n846,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1021, n1022, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1382, n1383, n1384, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147;
  wire   [9:0] genblk1_0__mac_s;
  wire   [9:0] genblk1_0__mac_biasesStored;
  wire   [9:0] genblk1_1__mac_s;
  wire   [9:0] genblk1_1__mac_biasesStored;
  wire   [9:0] genblk1_2__mac_s;
  wire   [9:0] genblk1_2__mac_biasesStored;
  wire   [9:0] genblk1_3__mac_s;
  wire   [9:0] genblk1_3__mac_biasesStored;
  wire   [9:0] genblk1_4__mac_s;
  wire   [9:0] genblk1_4__mac_biasesStored;
  wire   [9:0] genblk1_5__mac_s;
  wire   [9:0] genblk1_5__mac_biasesStored;
  wire   [9:0] genblk1_6__mac_s;
  wire   [9:0] genblk1_6__mac_biasesStored;
  wire   [9:0] genblk1_7__mac_s;
  wire   [9:0] genblk1_7__mac_biasesStored;
  wire   [9:0] genblk1_8__mac_s;
  wire   [9:0] genblk1_8__mac_biasesStored;
  wire   [9:0] genblk1_9__mac_s;
  wire   [9:0] genblk1_9__mac_biasesStored;

  DFFSRX4TS genblk1_0__mac_S_reg_1_ ( .D(genblk1_0__mac_s[1]), .CK(clk), .SN(
        n1), .RN(n2), .Q(sumOut[1]) );
  DFFSRX4TS genblk1_1__mac_S_reg_1_ ( .D(genblk1_1__mac_s[1]), .CK(clk), .SN(
        n13), .RN(n14), .Q(sumOut[11]) );
  DFFSRX4TS genblk1_3__mac_S_reg_1_ ( .D(genblk1_3__mac_s[1]), .CK(clk), .SN(
        n37), .RN(n38), .Q(sumOut[31]) );
  DFFSRX4TS genblk1_4__mac_S_reg_1_ ( .D(genblk1_4__mac_s[1]), .CK(clk), .SN(
        n49), .RN(n50), .Q(sumOut[41]) );
  DFFSRX4TS genblk1_5__mac_S_reg_1_ ( .D(genblk1_5__mac_s[1]), .CK(clk), .SN(
        n61), .RN(n62), .Q(sumOut[51]) );
  DFFSRX4TS genblk1_7__mac_S_reg_1_ ( .D(genblk1_7__mac_s[1]), .CK(clk), .SN(
        n85), .RN(n86), .Q(sumOut[71]) );
  DFFSRX4TS genblk1_0__mac_S_reg_2_ ( .D(genblk1_0__mac_s[2]), .CK(clk), .SN(
        n3), .RN(n4), .Q(sumOut[2]) );
  DFFSRX4TS genblk1_1__mac_S_reg_2_ ( .D(genblk1_1__mac_s[2]), .CK(clk), .SN(
        n15), .RN(n16), .Q(sumOut[12]) );
  DFFSRX4TS genblk1_1__mac_S_reg_3_ ( .D(genblk1_1__mac_s[3]), .CK(clk), .SN(
        n17), .RN(n18), .Q(sumOut[13]) );
  DFFSRX4TS genblk1_2__mac_S_reg_2_ ( .D(genblk1_2__mac_s[2]), .CK(clk), .SN(
        n27), .RN(n28), .Q(sumOut[22]) );
  DFFSRX4TS genblk1_2__mac_S_reg_3_ ( .D(genblk1_2__mac_s[3]), .CK(clk), .SN(
        n29), .RN(n30), .Q(sumOut[23]) );
  DFFSRX4TS genblk1_3__mac_S_reg_2_ ( .D(genblk1_3__mac_s[2]), .CK(clk), .SN(
        n39), .RN(n40), .Q(sumOut[32]) );
  DFFSRX4TS genblk1_3__mac_S_reg_3_ ( .D(genblk1_3__mac_s[3]), .CK(clk), .SN(
        n41), .RN(n42), .Q(sumOut[33]) );
  DFFSRX4TS genblk1_4__mac_S_reg_2_ ( .D(genblk1_4__mac_s[2]), .CK(clk), .SN(
        n51), .RN(n52), .Q(sumOut[42]) );
  DFFSRX4TS genblk1_4__mac_S_reg_3_ ( .D(genblk1_4__mac_s[3]), .CK(clk), .SN(
        n53), .RN(n54), .Q(sumOut[43]) );
  DFFSRX4TS genblk1_5__mac_S_reg_2_ ( .D(genblk1_5__mac_s[2]), .CK(clk), .SN(
        n63), .RN(n64), .Q(sumOut[52]) );
  DFFSRX4TS genblk1_5__mac_S_reg_3_ ( .D(genblk1_5__mac_s[3]), .CK(clk), .SN(
        n65), .RN(n66), .Q(sumOut[53]) );
  DFFSRX4TS genblk1_7__mac_S_reg_2_ ( .D(genblk1_7__mac_s[2]), .CK(clk), .SN(
        n87), .RN(n88), .Q(sumOut[72]) );
  DFFSRX4TS genblk1_7__mac_S_reg_3_ ( .D(genblk1_7__mac_s[3]), .CK(clk), .SN(
        n89), .RN(n90), .Q(sumOut[73]) );
  DFFSRX4TS genblk1_8__mac_S_reg_2_ ( .D(genblk1_8__mac_s[2]), .CK(clk), .SN(
        n99), .RN(n100), .Q(sumOut[82]) );
  DFFSRX4TS genblk1_8__mac_S_reg_3_ ( .D(genblk1_8__mac_s[3]), .CK(clk), .SN(
        n101), .RN(n102), .Q(sumOut[83]) );
  DFFSRX4TS genblk1_9__mac_S_reg_2_ ( .D(genblk1_9__mac_s[2]), .CK(clk), .SN(
        n111), .RN(n112), .Q(sumOut[92]) );
  DFFSRX4TS genblk1_9__mac_S_reg_3_ ( .D(genblk1_9__mac_s[3]), .CK(clk), .SN(
        n113), .RN(n114), .Q(sumOut[93]) );
  DFFSRX4TS genblk1_0__mac_S_reg_4_ ( .D(genblk1_0__mac_s[4]), .CK(clk), .SN(
        n7), .RN(n8), .Q(sumOut[4]), .QN(n462) );
  DFFSRX4TS genblk1_1__mac_S_reg_4_ ( .D(genblk1_1__mac_s[4]), .CK(clk), .SN(
        n19), .RN(n20), .Q(sumOut[14]) );
  DFFSRX4TS genblk1_2__mac_S_reg_4_ ( .D(genblk1_2__mac_s[4]), .CK(clk), .SN(
        n31), .RN(n32), .Q(sumOut[24]) );
  DFFSRX4TS genblk1_3__mac_S_reg_4_ ( .D(genblk1_3__mac_s[4]), .CK(clk), .SN(
        n43), .RN(n44), .Q(sumOut[34]) );
  DFFSRX4TS genblk1_4__mac_S_reg_4_ ( .D(genblk1_4__mac_s[4]), .CK(clk), .SN(
        n55), .RN(n56), .Q(sumOut[44]) );
  DFFSRX4TS genblk1_6__mac_S_reg_4_ ( .D(genblk1_6__mac_s[4]), .CK(clk), .SN(
        n79), .RN(n80), .Q(sumOut[64]) );
  DFFSRX4TS genblk1_7__mac_S_reg_4_ ( .D(genblk1_7__mac_s[4]), .CK(clk), .SN(
        n91), .RN(n92), .Q(sumOut[74]) );
  DFFSRX4TS genblk1_8__mac_S_reg_4_ ( .D(genblk1_8__mac_s[4]), .CK(clk), .SN(
        n103), .RN(n104), .Q(sumOut[84]) );
  DFFSRX4TS genblk1_9__mac_S_reg_4_ ( .D(genblk1_9__mac_s[4]), .CK(clk), .SN(
        n115), .RN(n116), .Q(sumOut[94]) );
  DFFSRX4TS genblk1_0__mac_S_reg_5_ ( .D(genblk1_0__mac_s[5]), .CK(clk), .SN(
        n532), .RN(n542), .Q(sumOut[5]) );
  DFFSRX4TS genblk1_2__mac_S_reg_5_ ( .D(genblk1_2__mac_s[5]), .CK(clk), .SN(
        n2131), .RN(n541), .Q(sumOut[25]), .QN(n457) );
  DFFSRX4TS genblk1_4__mac_S_reg_5_ ( .D(genblk1_4__mac_s[5]), .CK(clk), .SN(
        n528), .RN(n544), .Q(sumOut[45]), .QN(n456) );
  DFFSRX4TS genblk1_7__mac_S_reg_5_ ( .D(genblk1_7__mac_s[5]), .CK(clk), .SN(
        n524), .RN(n545), .Q(sumOut[75]) );
  DFFSRX4TS genblk1_9__mac_S_reg_5_ ( .D(genblk1_9__mac_s[5]), .CK(clk), .SN(
        n538), .RN(n118), .Q(sumOut[95]), .QN(n463) );
  DFFSRX4TS genblk1_0__mac_S_reg_6_ ( .D(genblk1_0__mac_s[6]), .CK(clk), .SN(
        n531), .RN(n542), .Q(sumOut[6]) );
  DFFSRX4TS genblk1_7__mac_S_reg_6_ ( .D(genblk1_7__mac_s[6]), .CK(clk), .SN(
        n523), .RN(n545), .Q(sumOut[76]), .QN(n459) );
  TLATXLTS genblk1_0__mac_biasesStored_reg_0_ ( .G(n2147), .D(biasesIn[0]), 
        .Q(genblk1_0__mac_biasesStored[0]) );
  TLATXLTS genblk1_0__mac_biasesStored_reg_1_ ( .G(n2147), .D(biasesIn[1]), 
        .Q(genblk1_0__mac_biasesStored[1]) );
  TLATXLTS genblk1_0__mac_biasesStored_reg_2_ ( .G(n2147), .D(biasesIn[2]), 
        .Q(genblk1_0__mac_biasesStored[2]) );
  TLATXLTS genblk1_0__mac_biasesStored_reg_3_ ( .G(n2147), .D(biasesIn[3]), 
        .Q(genblk1_0__mac_biasesStored[3]) );
  TLATXLTS genblk1_0__mac_biasesStored_reg_4_ ( .G(n2126), .D(biasesIn[4]), 
        .Q(genblk1_0__mac_biasesStored[4]) );
  TLATXLTS genblk1_0__mac_biasesStored_reg_9_ ( .G(n2133), .D(biasesIn[5]), 
        .Q(genblk1_0__mac_biasesStored[9]) );
  TLATXLTS genblk1_1__mac_biasesStored_reg_0_ ( .G(n2133), .D(biasesIn[6]), 
        .Q(genblk1_1__mac_biasesStored[0]) );
  TLATXLTS genblk1_1__mac_biasesStored_reg_1_ ( .G(n2133), .D(biasesIn[7]), 
        .Q(genblk1_1__mac_biasesStored[1]) );
  TLATXLTS genblk1_1__mac_biasesStored_reg_2_ ( .G(n2146), .D(biasesIn[8]), 
        .Q(genblk1_1__mac_biasesStored[2]) );
  TLATXLTS genblk1_1__mac_biasesStored_reg_3_ ( .G(n2146), .D(biasesIn[9]), 
        .Q(genblk1_1__mac_biasesStored[3]) );
  TLATXLTS genblk1_1__mac_biasesStored_reg_4_ ( .G(n2146), .D(biasesIn[10]), 
        .Q(genblk1_1__mac_biasesStored[4]) );
  TLATXLTS genblk1_1__mac_biasesStored_reg_9_ ( .G(n2146), .D(biasesIn[11]), 
        .Q(genblk1_1__mac_biasesStored[9]) );
  TLATXLTS genblk1_2__mac_biasesStored_reg_0_ ( .G(n2145), .D(biasesIn[12]), 
        .Q(genblk1_2__mac_biasesStored[0]) );
  TLATXLTS genblk1_2__mac_biasesStored_reg_1_ ( .G(n2145), .D(biasesIn[13]), 
        .Q(genblk1_2__mac_biasesStored[1]) );
  TLATXLTS genblk1_2__mac_biasesStored_reg_2_ ( .G(n2145), .D(biasesIn[14]), 
        .Q(genblk1_2__mac_biasesStored[2]) );
  TLATXLTS genblk1_2__mac_biasesStored_reg_3_ ( .G(n2145), .D(biasesIn[15]), 
        .Q(genblk1_2__mac_biasesStored[3]) );
  TLATXLTS genblk1_2__mac_biasesStored_reg_4_ ( .G(n2144), .D(biasesIn[16]), 
        .Q(genblk1_2__mac_biasesStored[4]) );
  TLATXLTS genblk1_2__mac_biasesStored_reg_9_ ( .G(n2144), .D(biasesIn[17]), 
        .Q(genblk1_2__mac_biasesStored[9]) );
  TLATXLTS genblk1_3__mac_biasesStored_reg_0_ ( .G(n2144), .D(biasesIn[18]), 
        .Q(genblk1_3__mac_biasesStored[0]) );
  TLATXLTS genblk1_3__mac_biasesStored_reg_1_ ( .G(n2144), .D(biasesIn[19]), 
        .Q(genblk1_3__mac_biasesStored[1]) );
  TLATXLTS genblk1_3__mac_biasesStored_reg_2_ ( .G(n2143), .D(biasesIn[20]), 
        .Q(genblk1_3__mac_biasesStored[2]) );
  TLATXLTS genblk1_3__mac_biasesStored_reg_3_ ( .G(n2143), .D(biasesIn[21]), 
        .Q(genblk1_3__mac_biasesStored[3]) );
  TLATXLTS genblk1_3__mac_biasesStored_reg_4_ ( .G(n2143), .D(biasesIn[22]), 
        .Q(genblk1_3__mac_biasesStored[4]) );
  TLATXLTS genblk1_3__mac_biasesStored_reg_9_ ( .G(n2143), .D(biasesIn[23]), 
        .Q(genblk1_3__mac_biasesStored[9]) );
  TLATXLTS genblk1_4__mac_biasesStored_reg_0_ ( .G(n2142), .D(biasesIn[24]), 
        .Q(genblk1_4__mac_biasesStored[0]) );
  TLATXLTS genblk1_4__mac_biasesStored_reg_1_ ( .G(n2142), .D(biasesIn[25]), 
        .Q(genblk1_4__mac_biasesStored[1]) );
  TLATXLTS genblk1_4__mac_biasesStored_reg_2_ ( .G(n2142), .D(biasesIn[26]), 
        .Q(genblk1_4__mac_biasesStored[2]) );
  TLATXLTS genblk1_4__mac_biasesStored_reg_3_ ( .G(n2142), .D(biasesIn[27]), 
        .Q(genblk1_4__mac_biasesStored[3]) );
  TLATXLTS genblk1_4__mac_biasesStored_reg_4_ ( .G(n2141), .D(biasesIn[28]), 
        .Q(genblk1_4__mac_biasesStored[4]) );
  TLATXLTS genblk1_4__mac_biasesStored_reg_9_ ( .G(n2141), .D(biasesIn[29]), 
        .Q(genblk1_4__mac_biasesStored[9]) );
  TLATXLTS genblk1_5__mac_biasesStored_reg_0_ ( .G(n2141), .D(biasesIn[30]), 
        .Q(genblk1_5__mac_biasesStored[0]) );
  TLATXLTS genblk1_5__mac_biasesStored_reg_1_ ( .G(n2141), .D(biasesIn[31]), 
        .Q(genblk1_5__mac_biasesStored[1]) );
  TLATXLTS genblk1_5__mac_biasesStored_reg_2_ ( .G(n2140), .D(biasesIn[32]), 
        .Q(genblk1_5__mac_biasesStored[2]) );
  TLATXLTS genblk1_5__mac_biasesStored_reg_3_ ( .G(n2140), .D(biasesIn[33]), 
        .Q(genblk1_5__mac_biasesStored[3]) );
  TLATXLTS genblk1_5__mac_biasesStored_reg_4_ ( .G(n2140), .D(biasesIn[34]), 
        .Q(genblk1_5__mac_biasesStored[4]) );
  TLATXLTS genblk1_5__mac_biasesStored_reg_9_ ( .G(n2140), .D(biasesIn[35]), 
        .Q(genblk1_5__mac_biasesStored[9]) );
  TLATXLTS genblk1_6__mac_biasesStored_reg_0_ ( .G(n2139), .D(biasesIn[36]), 
        .Q(genblk1_6__mac_biasesStored[0]) );
  TLATXLTS genblk1_6__mac_biasesStored_reg_1_ ( .G(n2139), .D(biasesIn[37]), 
        .Q(genblk1_6__mac_biasesStored[1]) );
  TLATXLTS genblk1_6__mac_biasesStored_reg_2_ ( .G(n2139), .D(biasesIn[38]), 
        .Q(genblk1_6__mac_biasesStored[2]) );
  TLATXLTS genblk1_6__mac_biasesStored_reg_3_ ( .G(n2139), .D(biasesIn[39]), 
        .Q(genblk1_6__mac_biasesStored[3]) );
  TLATXLTS genblk1_6__mac_biasesStored_reg_4_ ( .G(n2138), .D(biasesIn[40]), 
        .Q(genblk1_6__mac_biasesStored[4]) );
  TLATXLTS genblk1_6__mac_biasesStored_reg_9_ ( .G(n2138), .D(biasesIn[41]), 
        .Q(genblk1_6__mac_biasesStored[9]) );
  TLATXLTS genblk1_7__mac_biasesStored_reg_0_ ( .G(n2138), .D(biasesIn[42]), 
        .Q(genblk1_7__mac_biasesStored[0]) );
  TLATXLTS genblk1_7__mac_biasesStored_reg_1_ ( .G(n2138), .D(biasesIn[43]), 
        .Q(genblk1_7__mac_biasesStored[1]) );
  TLATXLTS genblk1_7__mac_biasesStored_reg_2_ ( .G(n2137), .D(biasesIn[44]), 
        .Q(genblk1_7__mac_biasesStored[2]) );
  TLATXLTS genblk1_7__mac_biasesStored_reg_3_ ( .G(n2137), .D(biasesIn[45]), 
        .Q(genblk1_7__mac_biasesStored[3]) );
  TLATXLTS genblk1_7__mac_biasesStored_reg_4_ ( .G(n2137), .D(biasesIn[46]), 
        .Q(genblk1_7__mac_biasesStored[4]) );
  TLATXLTS genblk1_7__mac_biasesStored_reg_9_ ( .G(n2137), .D(biasesIn[47]), 
        .Q(genblk1_7__mac_biasesStored[9]) );
  TLATXLTS genblk1_8__mac_biasesStored_reg_0_ ( .G(n2136), .D(biasesIn[48]), 
        .Q(genblk1_8__mac_biasesStored[0]) );
  TLATXLTS genblk1_8__mac_biasesStored_reg_1_ ( .G(n2136), .D(biasesIn[49]), 
        .Q(genblk1_8__mac_biasesStored[1]) );
  TLATXLTS genblk1_8__mac_biasesStored_reg_2_ ( .G(n2136), .D(biasesIn[50]), 
        .Q(genblk1_8__mac_biasesStored[2]) );
  TLATXLTS genblk1_8__mac_biasesStored_reg_3_ ( .G(n2136), .D(biasesIn[51]), 
        .Q(genblk1_8__mac_biasesStored[3]) );
  TLATXLTS genblk1_8__mac_biasesStored_reg_4_ ( .G(n2135), .D(biasesIn[52]), 
        .Q(genblk1_8__mac_biasesStored[4]) );
  TLATXLTS genblk1_8__mac_biasesStored_reg_9_ ( .G(n2135), .D(biasesIn[53]), 
        .Q(genblk1_8__mac_biasesStored[9]) );
  TLATXLTS genblk1_9__mac_biasesStored_reg_0_ ( .G(n2135), .D(biasesIn[54]), 
        .Q(genblk1_9__mac_biasesStored[0]) );
  TLATXLTS genblk1_9__mac_biasesStored_reg_1_ ( .G(n2135), .D(biasesIn[55]), 
        .Q(genblk1_9__mac_biasesStored[1]) );
  TLATXLTS genblk1_9__mac_biasesStored_reg_2_ ( .G(n2134), .D(biasesIn[56]), 
        .Q(genblk1_9__mac_biasesStored[2]) );
  TLATXLTS genblk1_9__mac_biasesStored_reg_3_ ( .G(n2134), .D(biasesIn[57]), 
        .Q(genblk1_9__mac_biasesStored[3]) );
  TLATXLTS genblk1_9__mac_biasesStored_reg_4_ ( .G(n2134), .D(biasesIn[58]), 
        .Q(genblk1_9__mac_biasesStored[4]) );
  TLATXLTS genblk1_9__mac_biasesStored_reg_9_ ( .G(n2134), .D(biasesIn[59]), 
        .Q(genblk1_9__mac_biasesStored[9]) );
  DFFSRX2TS genblk1_4__mac_S_reg_0_ ( .D(genblk1_4__mac_s[0]), .CK(clk), .SN(
        n59), .RN(n60), .Q(sumOut[40]) );
  DFFSRX2TS genblk1_5__mac_S_reg_0_ ( .D(genblk1_5__mac_s[0]), .CK(clk), .SN(
        n71), .RN(n72), .Q(sumOut[50]) );
  DFFSRX2TS genblk1_9__mac_S_reg_0_ ( .D(genblk1_9__mac_s[0]), .CK(clk), .SN(
        n119), .RN(n120), .Q(sumOut[90]) );
  DFFSRHQX4TS genblk1_9__mac_S_reg_7_ ( .D(genblk1_9__mac_s[7]), .CK(clk), 
        .SN(n538), .RN(n546), .Q(sumOut[97]) );
  DFFSRHQX4TS genblk1_9__mac_S_reg_8_ ( .D(genblk1_9__mac_s[8]), .CK(clk), 
        .SN(n538), .RN(n546), .Q(sumOut[98]) );
  DFFSRHQX4TS genblk1_3__mac_S_reg_9_ ( .D(genblk1_3__mac_s[9]), .CK(clk), 
        .SN(n530), .RN(n548), .Q(sumOut[39]) );
  DFFSRHQX4TS genblk1_1__mac_S_reg_8_ ( .D(genblk1_1__mac_s[8]), .CK(clk), 
        .SN(n533), .RN(n22), .Q(sumOut[18]) );
  DFFSRHQX4TS genblk1_1__mac_S_reg_7_ ( .D(genblk1_1__mac_s[7]), .CK(clk), 
        .SN(n534), .RN(n22), .Q(sumOut[17]) );
  DFFSRHQX4TS genblk1_3__mac_S_reg_8_ ( .D(genblk1_3__mac_s[8]), .CK(clk), 
        .SN(n530), .RN(n548), .Q(sumOut[38]) );
  DFFSRHQX4TS genblk1_4__mac_S_reg_8_ ( .D(genblk1_4__mac_s[8]), .CK(clk), 
        .SN(n529), .RN(n543), .Q(sumOut[48]) );
  DFFSRHQX4TS genblk1_9__mac_S_reg_9_ ( .D(genblk1_9__mac_s[9]), .CK(clk), 
        .SN(n538), .RN(n546), .Q(sumOut[99]) );
  DFFSRHQX4TS genblk1_4__mac_S_reg_9_ ( .D(genblk1_4__mac_s[9]), .CK(clk), 
        .SN(n529), .RN(n544), .Q(sumOut[49]) );
  DFFSRHQX4TS genblk1_4__mac_S_reg_7_ ( .D(genblk1_4__mac_s[7]), .CK(clk), 
        .SN(n529), .RN(n543), .Q(sumOut[47]) );
  DFFSRHQX4TS genblk1_6__mac_S_reg_2_ ( .D(genblk1_6__mac_s[2]), .CK(clk), 
        .SN(n75), .RN(n76), .Q(sumOut[62]) );
  DFFSRHQX4TS genblk1_6__mac_S_reg_5_ ( .D(genblk1_6__mac_s[5]), .CK(clk), 
        .SN(n525), .RN(n2132), .Q(sumOut[65]) );
  DFFSRHQX4TS genblk1_5__mac_S_reg_5_ ( .D(genblk1_5__mac_s[5]), .CK(clk), 
        .SN(n527), .RN(n547), .Q(sumOut[55]) );
  DFFSRHQX4TS genblk1_3__mac_S_reg_5_ ( .D(genblk1_3__mac_s[5]), .CK(clk), 
        .SN(n530), .RN(n549), .Q(sumOut[35]) );
  DFFSRHQX4TS genblk1_5__mac_S_reg_9_ ( .D(genblk1_5__mac_s[9]), .CK(clk), 
        .SN(n527), .RN(n547), .Q(sumOut[59]) );
  DFFSRHQX4TS genblk1_6__mac_S_reg_6_ ( .D(genblk1_6__mac_s[6]), .CK(clk), 
        .SN(n525), .RN(n82), .Q(sumOut[66]) );
  DFFSRHQX4TS genblk1_6__mac_S_reg_8_ ( .D(genblk1_6__mac_s[8]), .CK(clk), 
        .SN(n81), .RN(n2132), .Q(sumOut[68]) );
  DFFSRHQX4TS genblk1_1__mac_S_reg_5_ ( .D(genblk1_1__mac_s[5]), .CK(clk), 
        .SN(n534), .RN(n551), .Q(sumOut[15]) );
  DFFSRHQX4TS genblk1_6__mac_S_reg_7_ ( .D(genblk1_6__mac_s[7]), .CK(clk), 
        .SN(n81), .RN(n2132), .Q(sumOut[67]) );
  DFFSRHQX4TS genblk1_6__mac_S_reg_9_ ( .D(genblk1_6__mac_s[9]), .CK(clk), 
        .SN(n81), .RN(n2132), .Q(sumOut[69]) );
  DFFSRHQX4TS genblk1_7__mac_S_reg_8_ ( .D(genblk1_7__mac_s[8]), .CK(clk), 
        .SN(n524), .RN(n94), .Q(sumOut[78]) );
  DFFSRHQX4TS genblk1_0__mac_S_reg_9_ ( .D(genblk1_0__mac_s[9]), .CK(clk), 
        .SN(n532), .RN(n10), .Q(sumOut[9]) );
  DFFSRHQX4TS genblk1_8__mac_S_reg_8_ ( .D(genblk1_8__mac_s[8]), .CK(clk), 
        .SN(n536), .RN(n550), .Q(sumOut[88]) );
  DFFSRHQX4TS genblk1_1__mac_S_reg_9_ ( .D(genblk1_1__mac_s[9]), .CK(clk), 
        .SN(n534), .RN(n22), .Q(sumOut[19]) );
  DFFSRHQX4TS genblk1_1__mac_S_reg_6_ ( .D(genblk1_1__mac_s[6]), .CK(clk), 
        .SN(n534), .RN(n551), .Q(sumOut[16]) );
  DFFSRHQX4TS genblk1_7__mac_S_reg_9_ ( .D(genblk1_7__mac_s[9]), .CK(clk), 
        .SN(n524), .RN(n94), .Q(sumOut[79]) );
  DFFSRHQX4TS genblk1_3__mac_S_reg_7_ ( .D(genblk1_3__mac_s[7]), .CK(clk), 
        .SN(n45), .RN(n548), .Q(sumOut[37]) );
  DFFSRHQX4TS genblk1_5__mac_S_reg_8_ ( .D(genblk1_5__mac_s[8]), .CK(clk), 
        .SN(n527), .RN(n547), .Q(sumOut[58]) );
  DFFSRHQX4TS genblk1_2__mac_S_reg_8_ ( .D(genblk1_2__mac_s[8]), .CK(clk), 
        .SN(n2131), .RN(n541), .Q(sumOut[28]) );
  DFFSRHQX4TS genblk1_2__mac_S_reg_7_ ( .D(genblk1_2__mac_s[7]), .CK(clk), 
        .SN(n2131), .RN(n541), .Q(sumOut[27]) );
  DFFSRHQX4TS genblk1_5__mac_S_reg_7_ ( .D(genblk1_5__mac_s[7]), .CK(clk), 
        .SN(n527), .RN(n547), .Q(sumOut[57]) );
  DFFSRHQX4TS genblk1_0__mac_S_reg_7_ ( .D(genblk1_0__mac_s[7]), .CK(clk), 
        .SN(n532), .RN(n10), .Q(sumOut[7]) );
  DFFSRHQX4TS genblk1_0__mac_S_reg_8_ ( .D(genblk1_0__mac_s[8]), .CK(clk), 
        .SN(n532), .RN(n10), .Q(sumOut[8]) );
  DFFSRHQX4TS genblk1_7__mac_S_reg_7_ ( .D(genblk1_7__mac_s[7]), .CK(clk), 
        .SN(n524), .RN(n94), .Q(sumOut[77]) );
  DFFSRHQX4TS genblk1_2__mac_S_reg_9_ ( .D(genblk1_2__mac_s[9]), .CK(clk), 
        .SN(n2130), .RN(n541), .Q(sumOut[29]) );
  DFFSRHQX4TS genblk1_8__mac_S_reg_7_ ( .D(genblk1_8__mac_s[7]), .CK(clk), 
        .SN(n105), .RN(n106), .Q(sumOut[87]) );
  DFFSRHQX4TS genblk1_8__mac_S_reg_9_ ( .D(genblk1_8__mac_s[9]), .CK(clk), 
        .SN(n105), .RN(n106), .Q(sumOut[89]) );
  DFFSRHQX2TS genblk1_9__mac_S_reg_6_ ( .D(genblk1_9__mac_s[6]), .CK(clk), 
        .SN(n537), .RN(n118), .Q(sumOut[96]) );
  DFFSRHQX2TS genblk1_4__mac_S_reg_6_ ( .D(genblk1_4__mac_s[6]), .CK(clk), 
        .SN(n529), .RN(n543), .Q(sumOut[46]) );
  DFFSRHQX4TS genblk1_5__mac_S_reg_6_ ( .D(genblk1_5__mac_s[6]), .CK(clk), 
        .SN(n526), .RN(n70), .Q(sumOut[56]) );
  DFFSRX2TS genblk1_9__mac_S_reg_1_ ( .D(genblk1_9__mac_s[1]), .CK(clk), .SN(
        n109), .RN(n110), .Q(sumOut[91]) );
  DFFSRHQX2TS genblk1_8__mac_S_reg_0_ ( .D(genblk1_8__mac_s[0]), .CK(clk), 
        .SN(n107), .RN(n108), .Q(sumOut[80]) );
  DFFSRHQX2TS genblk1_1__mac_S_reg_0_ ( .D(genblk1_1__mac_s[0]), .CK(clk), 
        .SN(n23), .RN(n24), .Q(sumOut[10]) );
  DFFSRHQX2TS genblk1_8__mac_S_reg_5_ ( .D(genblk1_8__mac_s[5]), .CK(clk), 
        .SN(n536), .RN(n550), .Q(sumOut[85]) );
  DFFSRHQX2TS genblk1_3__mac_S_reg_6_ ( .D(genblk1_3__mac_s[6]), .CK(clk), 
        .SN(n530), .RN(n549), .Q(sumOut[36]) );
  DFFSRHQX2TS genblk1_8__mac_S_reg_6_ ( .D(genblk1_8__mac_s[6]), .CK(clk), 
        .SN(n105), .RN(n106), .Q(sumOut[86]) );
  DFFSRHQX2TS genblk1_2__mac_S_reg_6_ ( .D(genblk1_2__mac_s[6]), .CK(clk), 
        .SN(n2130), .RN(n540), .Q(sumOut[26]) );
  DFFSRX2TS genblk1_0__mac_S_reg_0_ ( .D(genblk1_0__mac_s[0]), .CK(clk), .SN(
        n11), .RN(n12), .Q(sumOut[0]) );
  DFFSRX2TS genblk1_6__mac_S_reg_0_ ( .D(genblk1_6__mac_s[0]), .CK(clk), .SN(
        n83), .RN(n84), .Q(sumOut[60]) );
  DFFSRX2TS genblk1_3__mac_S_reg_0_ ( .D(genblk1_3__mac_s[0]), .CK(clk), .SN(
        n47), .RN(n48), .Q(sumOut[30]) );
  DFFSRX2TS genblk1_2__mac_S_reg_0_ ( .D(genblk1_2__mac_s[0]), .CK(clk), .SN(
        n35), .RN(n36), .Q(sumOut[20]) );
  DFFSRX2TS genblk1_7__mac_S_reg_0_ ( .D(genblk1_7__mac_s[0]), .CK(clk), .SN(
        n95), .RN(n96), .Q(sumOut[70]) );
  DFFSRX2TS genblk1_6__mac_S_reg_1_ ( .D(genblk1_6__mac_s[1]), .CK(clk), .SN(
        n73), .RN(n74), .Q(sumOut[61]) );
  DFFSRX2TS genblk1_2__mac_S_reg_1_ ( .D(genblk1_2__mac_s[1]), .CK(clk), .SN(
        n25), .RN(n26), .Q(sumOut[21]) );
  DFFSRX2TS genblk1_8__mac_S_reg_1_ ( .D(genblk1_8__mac_s[1]), .CK(clk), .SN(
        n97), .RN(n98), .Q(sumOut[81]) );
  DFFSRX2TS genblk1_6__mac_S_reg_3_ ( .D(genblk1_6__mac_s[3]), .CK(clk), .SN(
        n77), .RN(n78), .Q(sumOut[63]) );
  DFFSRX2TS genblk1_0__mac_S_reg_3_ ( .D(genblk1_0__mac_s[3]), .CK(clk), .SN(
        n5), .RN(n6), .Q(sumOut[3]) );
  DFFSRX2TS genblk1_5__mac_S_reg_4_ ( .D(genblk1_5__mac_s[4]), .CK(clk), .SN(
        n67), .RN(n68), .Q(sumOut[54]) );
  CLKAND2X2TS U121 ( .A(n1847), .B(n1856), .Y(genblk1_1__mac_s[0]) );
  CLKAND2X2TS U122 ( .A(n1979), .B(n1977), .Y(n1722) );
  CLKAND2X2TS U123 ( .A(n1729), .B(n1728), .Y(n1730) );
  CLKAND2X2TS U124 ( .A(n1791), .B(n1789), .Y(n1785) );
  CLKAND2X2TS U125 ( .A(n1806), .B(n1805), .Y(n1807) );
  CLKAND2X2TS U126 ( .A(n269), .B(n1749), .Y(n1750) );
  CLKAND2X2TS U127 ( .A(n834), .B(n833), .Y(n835) );
  CLKBUFX2TS U128 ( .A(n1491), .Y(n1733) );
  INVX2TS U129 ( .A(n1158), .Y(n2075) );
  INVX1TS U130 ( .A(n2073), .Y(n181) );
  AOI21X2TS U131 ( .A0(n1407), .A1(n1406), .B0(n1405), .Y(n1408) );
  BUFX3TS U132 ( .A(n1560), .Y(n1457) );
  OR2X4TS U133 ( .A(n226), .B(sumOut[94]), .Y(n2073) );
  OAI21X2TS U134 ( .A0(n1848), .A1(n1851), .B0(n1850), .Y(n1489) );
  OR2X4TS U135 ( .A(n956), .B(n955), .Y(n1741) );
  OR2X4TS U136 ( .A(n1165), .B(n1164), .Y(n1525) );
  NAND2X4TS U137 ( .A(n159), .B(n158), .Y(n1832) );
  NAND2X1TS U138 ( .A(n659), .B(n658), .Y(n1884) );
  INVX2TS U139 ( .A(n1784), .Y(n1782) );
  NAND2X1TS U140 ( .A(n714), .B(sumOut[63]), .Y(n2000) );
  NOR2X1TS U141 ( .A(sumOut[79]), .B(n1515), .Y(n1514) );
  OAI2BB1X1TS U142 ( .A0N(n1836), .A1N(n1835), .B0(n310), .Y(n1837) );
  NOR2X4TS U143 ( .A(n1549), .B(n1548), .Y(n1708) );
  INVX1TS U144 ( .A(n1613), .Y(n158) );
  AOI21X2TS U145 ( .A0(n1901), .A1(n1899), .B0(n1361), .Y(n1915) );
  INVX3TS U146 ( .A(n1614), .Y(n159) );
  OAI21X1TS U147 ( .A0(n1835), .A1(n1836), .B0(sumOut[8]), .Y(n310) );
  OAI2BB1X2TS U148 ( .A0N(sumOut[55]), .A1N(n432), .B0(n828), .Y(n830) );
  OAI2BB1X2TS U149 ( .A0N(n906), .A1N(sumOut[15]), .B0(n861), .Y(n926) );
  OAI2BB1X2TS U150 ( .A0N(n148), .A1N(n1712), .B0(n164), .Y(n1721) );
  XOR2X2TS U151 ( .A(n1835), .B(n311), .Y(n1613) );
  XOR2X1TS U152 ( .A(n1797), .B(n1780), .Y(n1783) );
  OAI21X1TS U153 ( .A0(n1948), .A1(n1951), .B0(n1949), .Y(n1933) );
  NAND2X4TS U154 ( .A(n144), .B(n143), .Y(n1899) );
  INVX1TS U155 ( .A(n462), .Y(n171) );
  NOR2X2TS U156 ( .A(sumOut[11]), .B(n913), .Y(n1853) );
  NOR2X1TS U157 ( .A(sumOut[31]), .B(n1356), .Y(n1917) );
  NAND2X1TS U158 ( .A(sumOut[82]), .B(n1661), .Y(n2038) );
  NAND2X1TS U159 ( .A(sumOut[2]), .B(n1448), .Y(n1809) );
  NAND2X1TS U160 ( .A(sumOut[20]), .B(n1867), .Y(n1877) );
  CLKINVX2TS U161 ( .A(n1332), .Y(n1335) );
  OAI21X2TS U162 ( .A0(n753), .A1(n754), .B0(sumOut[66]), .Y(n752) );
  OAI21X2TS U163 ( .A0(n1753), .A1(n1754), .B0(sumOut[86]), .Y(n1752) );
  OAI21X2TS U164 ( .A0(n1586), .A1(n1585), .B0(sumOut[6]), .Y(n1584) );
  NAND2X1TS U165 ( .A(sumOut[60]), .B(n1994), .Y(n2007) );
  OAI21X1TS U166 ( .A0(sumOut[45]), .A1(n1034), .B0(n1036), .Y(n972) );
  NAND2X1TS U167 ( .A(sumOut[10]), .B(n1846), .Y(n1856) );
  OAI2BB1X1TS U168 ( .A0N(n463), .A1N(n1116), .B0(n1115), .Y(n1117) );
  OAI21X1TS U169 ( .A0(n1003), .A1(n1002), .B0(sumOut[47]), .Y(n1004) );
  XOR2X2TS U170 ( .A(n428), .B(n1450), .Y(n1453) );
  CLKINVX1TS U171 ( .A(sumOut[93]), .Y(n131) );
  NAND2X1TS U172 ( .A(sumOut[70]), .B(n2020), .Y(n2036) );
  OAI21X2TS U173 ( .A0(sumOut[55]), .A1(n432), .B0(n827), .Y(n828) );
  XOR2X1TS U174 ( .A(n1836), .B(sumOut[8]), .Y(n311) );
  OAI2BB1X4TS U175 ( .A0N(n1359), .A1N(n1358), .B0(n361), .Y(n1373) );
  XOR2X1TS U176 ( .A(n1798), .B(sumOut[88]), .Y(n1780) );
  XOR2X1TS U177 ( .A(n1892), .B(sumOut[28]), .Y(n657) );
  NAND2X4TS U178 ( .A(n2067), .B(n2069), .Y(n354) );
  CLKINVX1TS U179 ( .A(sumOut[32]), .Y(n143) );
  OR2X1TS U180 ( .A(n245), .B(n1714), .Y(n1985) );
  INVX4TS U181 ( .A(n1360), .Y(n144) );
  NAND2X1TS U182 ( .A(sumOut[11]), .B(n913), .Y(n1854) );
  BUFX6TS U183 ( .A(n1640), .Y(n1674) );
  BUFX2TS U184 ( .A(n1697), .Y(n1700) );
  NOR2X1TS U185 ( .A(n678), .B(n1180), .Y(n2020) );
  OAI2BB1X1TS U186 ( .A0N(n1639), .A1N(n1629), .B0(n1638), .Y(n1673) );
  NAND2X4TS U187 ( .A(n426), .B(n335), .Y(n1380) );
  OAI2BB1X2TS U188 ( .A0N(n1137), .A1N(n1136), .B0(n1135), .Y(n1141) );
  NAND2X4TS U189 ( .A(n185), .B(n186), .Y(n1332) );
  INVX2TS U190 ( .A(n1232), .Y(n431) );
  CLKBUFX2TS U191 ( .A(sumOut[46]), .Y(n977) );
  CLKBUFX2TS U192 ( .A(n826), .Y(n432) );
  BUFX3TS U193 ( .A(n1713), .Y(n148) );
  OR2X2TS U194 ( .A(n1715), .B(n656), .Y(n1892) );
  XNOR2X1TS U195 ( .A(n912), .B(n328), .Y(n913) );
  XOR2X1TS U196 ( .A(n702), .B(n701), .Y(n704) );
  XOR2X2TS U197 ( .A(n1226), .B(n1225), .Y(n1227) );
  ADDFHX2TS U198 ( .A(n1612), .B(n1611), .CI(n1610), .CO(n1835), .S(n1607) );
  ADDFHX2TS U199 ( .A(n1395), .B(n1394), .CI(n1393), .CO(n1410), .S(n1398) );
  CLKINVX1TS U200 ( .A(sumOut[27]), .Y(n153) );
  NAND3X2TS U201 ( .A(n175), .B(n174), .C(n176), .Y(n1039) );
  OR2X1TS U202 ( .A(n245), .B(n1499), .Y(n1512) );
  CLKBUFX2TS U203 ( .A(n579), .Y(n413) );
  CLKBUFX3TS U204 ( .A(n1214), .Y(n1051) );
  INVX2TS U205 ( .A(n707), .Y(n708) );
  OAI2BB1X2TS U206 ( .A0N(n1244), .A1N(n1243), .B0(n1242), .Y(n1248) );
  NAND2X1TS U207 ( .A(sumOut[90]), .B(n2070), .Y(n2083) );
  OAI21X2TS U208 ( .A0(n1758), .A1(n1757), .B0(n1755), .Y(n1756) );
  CLKBUFX2TS U209 ( .A(n502), .Y(n207) );
  XOR2X2TS U210 ( .A(n500), .B(n503), .Y(n481) );
  OAI21X2TS U211 ( .A0(n976), .A1(n975), .B0(n973), .Y(n974) );
  NAND2X4TS U212 ( .A(n324), .B(n1366), .Y(n426) );
  XOR2X2TS U213 ( .A(n1358), .B(n1359), .Y(n360) );
  NAND2X1TS U214 ( .A(n1246), .B(n1245), .Y(n1247) );
  NAND2X2TS U215 ( .A(n170), .B(n1025), .Y(n176) );
  OR2X2TS U216 ( .A(n842), .B(n951), .Y(n953) );
  INVX1TS U217 ( .A(n284), .Y(n285) );
  INVX1TS U218 ( .A(n151), .Y(n1204) );
  NAND2X1TS U219 ( .A(n1338), .B(n1339), .Y(n320) );
  NOR2X1TS U220 ( .A(n596), .B(n557), .Y(n599) );
  NOR2X2TS U221 ( .A(n842), .B(n1124), .Y(n1137) );
  AND2X6TS U222 ( .A(n1021), .B(n1022), .Y(n1014) );
  INVX2TS U223 ( .A(n1245), .Y(n1243) );
  OAI2BB1X2TS U224 ( .A0N(n1447), .A1N(n1446), .B0(n377), .Y(n1452) );
  OAI2BB1X2TS U225 ( .A0N(n785), .A1N(n786), .B0(n784), .Y(n393) );
  CLKINVX2TS U226 ( .A(n1246), .Y(n1244) );
  CLKINVX2TS U227 ( .A(n1573), .Y(n1467) );
  OAI21X2TS U228 ( .A0(n865), .A1(n862), .B0(n863), .Y(n864) );
  NAND2X2TS U229 ( .A(n627), .B(n625), .Y(n453) );
  INVX2TS U230 ( .A(n512), .Y(n318) );
  NAND2BX2TS U231 ( .AN(n1124), .B(n1123), .Y(n1142) );
  NOR2X4TS U232 ( .A(n242), .B(n1689), .Y(n1758) );
  NAND2X1TS U233 ( .A(n627), .B(n626), .Y(n454) );
  NAND2X1TS U234 ( .A(n557), .B(n596), .Y(n597) );
  OR2X2TS U235 ( .A(n1659), .B(n1007), .Y(n975) );
  OR2X4TS U236 ( .A(n1443), .B(n878), .Y(n858) );
  CLKBUFX2TS U237 ( .A(n1026), .Y(n170) );
  OAI21X2TS U238 ( .A0(n1595), .A1(n1594), .B0(n1592), .Y(n1593) );
  XOR2X2TS U239 ( .A(n476), .B(n475), .Y(n317) );
  CLKBUFX2TS U240 ( .A(n696), .Y(n284) );
  XOR2X1TS U241 ( .A(n471), .B(n470), .Y(n468) );
  INVX1TS U242 ( .A(n276), .Y(n124) );
  OAI21X1TS U243 ( .A0(n1760), .A1(n167), .B0(n1761), .Y(n165) );
  NOR2X2TS U244 ( .A(n745), .B(n1205), .Y(n1201) );
  INVX2TS U245 ( .A(n1589), .Y(n156) );
  CLKINVX1TS U246 ( .A(n1543), .Y(n162) );
  XOR2X2TS U247 ( .A(n674), .B(n675), .Y(n697) );
  NOR2X2TS U248 ( .A(n842), .B(n990), .Y(n996) );
  NOR2X4TS U249 ( .A(n1591), .B(n383), .Y(n1589) );
  INVX4TS U250 ( .A(n1127), .Y(n1145) );
  OAI2BB1X2TS U251 ( .A0N(n822), .A1N(n821), .B0(n820), .Y(n1542) );
  AND2X2TS U252 ( .A(n605), .B(n606), .Y(n613) );
  OAI2BB1X2TS U253 ( .A0N(n424), .A1N(n363), .B0(n686), .Y(n687) );
  AND2X4TS U254 ( .A(n677), .B(n676), .Y(n672) );
  BUFX4TS U255 ( .A(n1344), .Y(n301) );
  INVX2TS U256 ( .A(n1323), .Y(n1343) );
  INVX4TS U257 ( .A(n1123), .Y(n1715) );
  NOR2X2TS U258 ( .A(n593), .B(n196), .Y(n591) );
  OAI21X2TS U259 ( .A0(n168), .A1(n850), .B0(n846), .Y(n849) );
  INVX1TS U260 ( .A(n1320), .Y(n313) );
  OAI21X1TS U261 ( .A0(n1107), .A1(n1106), .B0(n1104), .Y(n1105) );
  CLKBUFX2TS U262 ( .A(n611), .Y(n125) );
  OAI21X2TS U263 ( .A0(n732), .A1(n733), .B0(n357), .Y(n731) );
  NOR2X4TS U264 ( .A(n1618), .B(n889), .Y(n893) );
  OR2X2TS U265 ( .A(n188), .B(n951), .Y(n729) );
  AND2X4TS U266 ( .A(n1631), .B(n1632), .Y(n458) );
  AND2X4TS U267 ( .A(n900), .B(n899), .Y(n896) );
  NOR2X4TS U268 ( .A(n1692), .B(n1693), .Y(n1760) );
  NOR2X4TS U269 ( .A(n1625), .B(n1346), .Y(n1369) );
  NAND2X4TS U270 ( .A(n1329), .B(n981), .Y(n986) );
  OAI21X2TS U271 ( .A0(n915), .A1(n916), .B0(n914), .Y(n302) );
  NOR2X2TS U272 ( .A(n1633), .B(n604), .Y(n615) );
  NOR2X8TS U273 ( .A(n1207), .B(n1029), .Y(n1021) );
  NOR2X4TS U274 ( .A(n383), .B(n691), .Y(n693) );
  AND2X6TS U275 ( .A(n1691), .B(n282), .Y(n274) );
  NOR2X2TS U276 ( .A(n1434), .B(n1029), .Y(n1044) );
  NAND2X6TS U277 ( .A(n1695), .B(n1470), .Y(n1578) );
  NOR2X4TS U278 ( .A(n1214), .B(n823), .Y(n771) );
  INVX2TS U279 ( .A(n386), .Y(n1631) );
  INVX2TS U280 ( .A(n1125), .Y(n1128) );
  NOR2X4TS U281 ( .A(n1016), .B(n1421), .Y(n1575) );
  OR2X2TS U282 ( .A(n898), .B(n1327), .Y(n1321) );
  OR2X2TS U283 ( .A(n239), .B(n1150), .Y(n1102) );
  NOR2X2TS U284 ( .A(n1302), .B(n691), .Y(n675) );
  BUFX3TS U285 ( .A(n730), .Y(n357) );
  BUFX3TS U286 ( .A(n356), .Y(n135) );
  INVX6TS U287 ( .A(n1338), .Y(n276) );
  AND2X4TS U288 ( .A(n702), .B(n701), .Y(n707) );
  NAND2X4TS U289 ( .A(n264), .B(n146), .Y(n145) );
  NAND2X1TS U290 ( .A(n192), .B(n1018), .Y(n1027) );
  AND2X4TS U291 ( .A(n912), .B(n327), .Y(n914) );
  AND2X4TS U292 ( .A(n1691), .B(n1622), .Y(n1761) );
  AND2X4TS U293 ( .A(n1349), .B(n1350), .Y(n1364) );
  AND2X4TS U294 ( .A(n969), .B(n248), .Y(n598) );
  OR2X4TS U295 ( .A(n1207), .B(n243), .Y(n1685) );
  AND2X6TS U296 ( .A(n471), .B(n470), .Y(n474) );
  INVX2TS U297 ( .A(n781), .Y(n786) );
  INVX3TS U298 ( .A(n488), .Y(n512) );
  NAND2X4TS U299 ( .A(n203), .B(n959), .Y(n963) );
  NOR2X6TS U300 ( .A(n1432), .B(n1017), .Y(n966) );
  NAND2X4TS U301 ( .A(n388), .B(n338), .Y(n389) );
  NOR2X6TS U302 ( .A(n1619), .B(n886), .Y(n855) );
  NAND2X2TS U303 ( .A(n1109), .B(n1695), .Y(n1104) );
  NOR2X2TS U304 ( .A(n1434), .B(n601), .Y(n606) );
  AND2X4TS U305 ( .A(n189), .B(n851), .Y(n854) );
  NOR2X4TS U306 ( .A(n244), .B(n567), .Y(n626) );
  NOR2X4TS U307 ( .A(n1443), .B(n1692), .Y(n1629) );
  NOR2X4TS U308 ( .A(n1633), .B(n593), .Y(n574) );
  NOR2X2TS U309 ( .A(n1214), .B(n775), .Y(n802) );
  NOR2X2TS U310 ( .A(n1646), .B(n1633), .Y(n1634) );
  INVX6TS U311 ( .A(n202), .Y(n1625) );
  BUFX6TS U312 ( .A(n508), .Y(n338) );
  BUFX6TS U313 ( .A(n465), .Y(n1443) );
  INVX2TS U314 ( .A(n1195), .Y(n1186) );
  INVX2TS U315 ( .A(n662), .Y(n734) );
  INVX2TS U316 ( .A(n328), .Y(n327) );
  NOR2X2TS U317 ( .A(n1633), .B(n467), .Y(n470) );
  NOR2X2TS U318 ( .A(n1417), .B(n469), .Y(n471) );
  NAND2X4TS U319 ( .A(n767), .B(n193), .Y(n781) );
  AND2X4TS U320 ( .A(n491), .B(n767), .Y(n461) );
  INVX4TS U321 ( .A(n141), .Y(n1350) );
  NOR2X6TS U322 ( .A(n765), .B(n1340), .Y(n455) );
  NOR2X6TS U323 ( .A(n745), .B(n823), .Y(n822) );
  NOR2X2TS U324 ( .A(n1050), .B(n1207), .Y(n1049) );
  INVX2TS U325 ( .A(n241), .Y(n1622) );
  NAND2X6TS U326 ( .A(n991), .B(n853), .Y(n848) );
  INVX4TS U327 ( .A(n363), .Y(n688) );
  AND2X4TS U328 ( .A(n195), .B(n1426), .Y(n1430) );
  BUFX3TS U329 ( .A(n509), .Y(n388) );
  CLKBUFX2TS U330 ( .A(weightsIn[28]), .Y(n968) );
  NAND2X4TS U331 ( .A(n837), .B(n1469), .Y(n350) );
  NOR2X1TS U332 ( .A(n898), .B(n776), .Y(n807) );
  INVX2TS U333 ( .A(n282), .Y(n601) );
  INVX4TS U334 ( .A(n308), .Y(n307) );
  NAND2X2TS U335 ( .A(n200), .B(n1313), .Y(n375) );
  INVX2TS U336 ( .A(n139), .Y(n138) );
  INVX2TS U337 ( .A(n843), .Y(n853) );
  CLKINVX3TS U338 ( .A(n1322), .Y(n1324) );
  NAND2X2TS U339 ( .A(n1422), .B(n1691), .Y(n308) );
  AND2X4TS U340 ( .A(n211), .B(n263), .Y(n1307) );
  NAND2X2TS U341 ( .A(n837), .B(n200), .Y(n328) );
  NOR2X6TS U342 ( .A(n1432), .B(n1442), .Y(n139) );
  CLKBUFX2TS U343 ( .A(weightsIn[58]), .Y(n1109) );
  BUFX8TS U344 ( .A(n1340), .Y(n134) );
  NAND2X4TS U345 ( .A(n198), .B(n1426), .Y(n342) );
  INVX2TS U346 ( .A(n1030), .Y(n959) );
  NAND2X6TS U347 ( .A(n1251), .B(n489), .Y(n509) );
  INVX2TS U348 ( .A(n240), .Y(n241) );
  INVX2TS U349 ( .A(n887), .Y(n901) );
  NAND2X4TS U350 ( .A(n1469), .B(n1249), .Y(n356) );
  INVX2TS U351 ( .A(n337), .Y(n1308) );
  CLKBUFX2TS U352 ( .A(n1626), .Y(n364) );
  NAND2X4TS U353 ( .A(n1019), .B(n251), .Y(n141) );
  NAND2X4TS U354 ( .A(n491), .B(n1110), .Y(n508) );
  INVX6TS U355 ( .A(n189), .Y(n465) );
  INVX8TS U356 ( .A(n1469), .Y(n1432) );
  INVX2TS U357 ( .A(n1425), .Y(n1442) );
  BUFX8TS U358 ( .A(n190), .Y(n200) );
  BUFX3TS U359 ( .A(weightsIn[1]), .Y(n1426) );
  INVX2TS U360 ( .A(n1312), .Y(n1313) );
  BUFX3TS U361 ( .A(weightsIn[55]), .Y(n489) );
  INVX8TS U362 ( .A(n195), .Y(n196) );
  CLKBUFX2TS U363 ( .A(weightsIn[32]), .Y(n761) );
  INVX2TS U364 ( .A(n667), .Y(n662) );
  CLKBUFX2TS U365 ( .A(weightsIn[15]), .Y(n555) );
  CLKBUFX2TS U366 ( .A(weightsIn[57]), .Y(n1110) );
  INVX3TS U367 ( .A(n259), .Y(n260) );
  BUFX6TS U368 ( .A(n571), .Y(n969) );
  CLKBUFX2TS U369 ( .A(weightsIn[0]), .Y(n1425) );
  INVX2TS U370 ( .A(weightsIn[54]), .Y(n259) );
  INVX2TS U371 ( .A(weightsIn[52]), .Y(n1690) );
  INVX2TS U372 ( .A(weightsIn[37]), .Y(n256) );
  OAI2BB1X2TS U373 ( .A0N(n671), .A1N(n670), .B0(n669), .Y(n715) );
  OAI21X2TS U374 ( .A0(n502), .A1(n503), .B0(n500), .Y(n501) );
  NAND2X1TS U375 ( .A(n2058), .B(n2046), .Y(n2047) );
  CLKINVX3TS U376 ( .A(n351), .Y(n397) );
  OAI2BB1X2TS U377 ( .A0N(n1450), .A1N(n428), .B0(n1435), .Y(n1473) );
  OAI21X4TS U378 ( .A0(n1688), .A1(n1687), .B0(n1685), .Y(n1686) );
  INVX2TS U379 ( .A(n1264), .Y(n420) );
  XOR2X1TS U380 ( .A(n1767), .B(n1766), .Y(genblk1_8__mac_s[7]) );
  INVX6TS U381 ( .A(n1108), .Y(n1303) );
  NAND2X2TS U382 ( .A(n2073), .B(n2072), .Y(n2074) );
  NAND2X4TS U383 ( .A(n711), .B(n710), .Y(n1991) );
  OAI21X2TS U384 ( .A0(n1970), .A1(n405), .B0(n411), .Y(n1975) );
  NOR2X2TS U385 ( .A(n480), .B(n479), .Y(n496) );
  NAND2X2TS U386 ( .A(n206), .B(n1997), .Y(n1998) );
  INVX8TS U387 ( .A(n200), .Y(n244) );
  XNOR2X1TS U388 ( .A(n126), .B(n128), .Y(genblk1_9__mac_s[8]) );
  OAI21X2TS U389 ( .A0(n1523), .A1(n2087), .B0(n1522), .Y(n126) );
  OAI21X2TS U390 ( .A0(n670), .A1(n671), .B0(n672), .Y(n669) );
  XOR2X1TS U391 ( .A(n1786), .B(n1785), .Y(genblk1_8__mac_s[8]) );
  OAI21X2TS U392 ( .A0(n1772), .A1(n1794), .B0(n1771), .Y(n1786) );
  XOR2X4TS U393 ( .A(n910), .B(n909), .Y(n295) );
  INVX8TS U394 ( .A(n1689), .Y(n370) );
  OAI2BB1X2TS U395 ( .A0N(n1217), .A1N(n1218), .B0(n1198), .Y(n1234) );
  INVX6TS U396 ( .A(n1196), .Y(n571) );
  XOR2X1TS U397 ( .A(n1551), .B(n1550), .Y(genblk1_5__mac_s[7]) );
  XOR2X1TS U398 ( .A(n1808), .B(n1807), .Y(genblk1_3__mac_s[7]) );
  XOR2X1TS U399 ( .A(n1731), .B(n1730), .Y(genblk1_7__mac_s[8]) );
  OAI21X1TS U400 ( .A0(n1727), .A1(n2024), .B0(n1726), .Y(n1731) );
  NAND2X2TS U401 ( .A(n353), .B(n1880), .Y(n1881) );
  XOR2X1TS U402 ( .A(n288), .B(n1989), .Y(genblk1_5__mac_s[9]) );
  OAI21X2TS U403 ( .A0(n1589), .A1(n1590), .B0(n1587), .Y(n1588) );
  INVX2TS U404 ( .A(n1683), .Y(n1681) );
  NAND2X4TS U405 ( .A(n194), .B(n1621), .Y(n351) );
  INVX8TS U406 ( .A(n490), .Y(n1108) );
  CLKINVX6TS U407 ( .A(n304), .Y(n1466) );
  OAI21X2TS U408 ( .A0(n1576), .A1(n1575), .B0(n1578), .Y(n1574) );
  NAND2X2TS U409 ( .A(n1403), .B(n1406), .Y(n1409) );
  INVX2TS U410 ( .A(n1403), .Y(n1392) );
  NOR2BX2TS U411 ( .AN(n1706), .B(n1708), .Y(n1550) );
  NOR2X4TS U412 ( .A(n594), .B(n1312), .Y(n1395) );
  OAI21X2TS U413 ( .A0(n445), .A1(n1380), .B0(n1378), .Y(n1379) );
  AND2X4TS U414 ( .A(n1354), .B(n1355), .Y(n1357) );
  OAI21X2TS U415 ( .A0(n1358), .A1(n1359), .B0(n1357), .Y(n361) );
  INVX2TS U416 ( .A(n199), .Y(n1651) );
  AND2X4TS U417 ( .A(n675), .B(n674), .Y(n696) );
  XOR2X4TS U418 ( .A(n822), .B(n819), .Y(n133) );
  BUFX20TS U419 ( .A(n760), .Y(n198) );
  INVX6TS U420 ( .A(n339), .Y(n1251) );
  NAND2X6TS U421 ( .A(n193), .B(n282), .Y(n334) );
  BUFX3TS U422 ( .A(n2022), .Y(n121) );
  NAND2X4TS U423 ( .A(n194), .B(n1250), .Y(n333) );
  CLKINVX6TS U424 ( .A(n888), .Y(n895) );
  OAI2BB1X4TS U425 ( .A0N(n910), .A1N(n909), .B0(n902), .Y(n446) );
  OAI21X4TS U426 ( .A0(n910), .A1(n909), .B0(n911), .Y(n902) );
  XOR2X4TS U427 ( .A(n860), .B(n444), .Y(n907) );
  AOI21X4TS U428 ( .A0(n1831), .A1(n1832), .B0(n1830), .Y(n136) );
  OAI21X4TS U429 ( .A0(n1815), .A1(n1603), .B0(n1602), .Y(n1831) );
  INVX12TS U430 ( .A(n877), .Y(n1016) );
  AND2X8TS U431 ( .A(n877), .B(weightsIn[24]), .Y(n1026) );
  BUFX4TS U432 ( .A(n516), .Y(n316) );
  XOR2X4TS U433 ( .A(n508), .B(n509), .Y(n494) );
  XOR2X4TS U434 ( .A(n122), .B(n980), .Y(n973) );
  XOR2X4TS U435 ( .A(n979), .B(n985), .Y(n122) );
  OAI21X4TS U436 ( .A0(n1286), .A1(n1078), .B0(n1079), .Y(n1091) );
  NOR2X8TS U437 ( .A(n1063), .B(n1062), .Y(n1078) );
  XOR2X4TS U438 ( .A(n992), .B(n1008), .Y(n1002) );
  OAI2BB1X4TS U439 ( .A0N(n988), .A1N(n989), .B0(n987), .Y(n1008) );
  INVX8TS U440 ( .A(n571), .Y(n1302) );
  INVX16TS U441 ( .A(n1302), .Y(n1691) );
  INVX6TS U442 ( .A(n1196), .Y(n490) );
  BUFX12TS U443 ( .A(n490), .Y(n1469) );
  CLKINVX1TS U444 ( .A(n123), .Y(n883) );
  XNOR2X4TS U445 ( .A(n123), .B(n882), .Y(n885) );
  NAND2X4TS U446 ( .A(n149), .B(n893), .Y(n123) );
  XNOR2X4TS U447 ( .A(n998), .B(n1003), .Y(n1063) );
  NOR2X4TS U448 ( .A(n1388), .B(n1387), .Y(n1904) );
  INVX8TS U449 ( .A(n877), .Y(n1262) );
  NOR2X6TS U450 ( .A(n1017), .B(n1262), .Y(n988) );
  NAND2X4TS U451 ( .A(n194), .B(n1311), .Y(n1322) );
  INVX6TS U452 ( .A(n1108), .Y(n491) );
  XOR2X4TS U453 ( .A(n1339), .B(n276), .Y(n1330) );
  NOR2X8TS U454 ( .A(n134), .B(n1312), .Y(n1338) );
  NOR2X6TS U455 ( .A(n1923), .B(n1925), .Y(n1386) );
  NOR2X8TS U456 ( .A(n1383), .B(n1384), .Y(n1925) );
  OAI21X4TS U457 ( .A0(n1324), .A1(n1325), .B0(n1323), .Y(n382) );
  OAI21X2TS U458 ( .A0(n1339), .A1(n124), .B0(n1337), .Y(n321) );
  INVX4TS U459 ( .A(n1365), .Y(n324) );
  NOR2X6TS U460 ( .A(n1637), .B(sumOut[84]), .Y(n2059) );
  INVX4TS U461 ( .A(n1196), .Y(n760) );
  NOR2X8TS U462 ( .A(n1418), .B(n886), .Y(n865) );
  INVX6TS U463 ( .A(n1347), .Y(n1618) );
  INVX12TS U464 ( .A(n1347), .Y(n1468) );
  INVX4TS U465 ( .A(layer2In[1]), .Y(n1196) );
  NOR2X4TS U466 ( .A(n1301), .B(n1302), .Y(n1349) );
  XOR2X4TS U467 ( .A(n1354), .B(n1355), .Y(n1356) );
  XOR2X1TS U468 ( .A(n1533), .B(n1532), .Y(genblk1_9__mac_s[7]) );
  XOR2X1TS U469 ( .A(n1176), .B(n1175), .Y(genblk1_9__mac_s[9]) );
  OAI21X4TS U470 ( .A0(n1155), .A1(n1156), .B0(n1154), .Y(n1157) );
  NOR2X8TS U471 ( .A(n518), .B(n519), .Y(n1155) );
  OAI21X2TS U472 ( .A0(n1983), .A1(n1982), .B0(n1981), .Y(n288) );
  INVX6TS U473 ( .A(n1108), .Y(n211) );
  NAND2X6TS U474 ( .A(n211), .B(n489), .Y(n479) );
  OAI2BB1X4TS U475 ( .A0N(n1543), .A1N(n1542), .B0(n294), .Y(n1712) );
  OAI21X4TS U476 ( .A0(n822), .A1(n821), .B0(n1535), .Y(n820) );
  INVX6TS U477 ( .A(n339), .Y(n194) );
  AOI21X4TS U478 ( .A0(n1386), .A1(n1909), .B0(n127), .Y(n1907) );
  OAI21X4TS U479 ( .A0(n1925), .A1(n1922), .B0(n1927), .Y(n127) );
  NAND2X1TS U480 ( .A(n1525), .B(n1524), .Y(n128) );
  INVX6TS U481 ( .A(n877), .Y(n1418) );
  CLKINVX6TS U482 ( .A(n333), .Y(n329) );
  OAI2BB1X2TS U483 ( .A0N(n1141), .A1N(n1140), .B0(n1139), .Y(n1165) );
  OAI21X2TS U484 ( .A0(n1006), .A1(n1005), .B0(n1004), .Y(n1065) );
  INVX8TS U485 ( .A(n592), .Y(n1310) );
  INVX8TS U486 ( .A(n1310), .Y(n202) );
  CLKINVX6TS U487 ( .A(n299), .Y(n298) );
  INVX8TS U488 ( .A(n1310), .Y(n203) );
  OAI2BB1X4TS U489 ( .A0N(n517), .A1N(n316), .B0(n129), .Y(n518) );
  OAI21X4TS U490 ( .A0(n316), .A1(n517), .B0(n514), .Y(n129) );
  BUFX16TS U491 ( .A(n592), .Y(n193) );
  CLKINVX3TS U492 ( .A(n770), .Y(n769) );
  XOR2X4TS U493 ( .A(n782), .B(n781), .Y(n763) );
  OAI21X4TS U494 ( .A0(n476), .A1(n475), .B0(n474), .Y(n478) );
  BUFX3TS U495 ( .A(n1707), .Y(n130) );
  INVX4TS U496 ( .A(n484), .Y(n132) );
  NAND2X4TS U497 ( .A(n132), .B(n131), .Y(n482) );
  XNOR2X4TS U498 ( .A(n133), .B(n1535), .Y(n817) );
  NAND2X4TS U499 ( .A(n307), .B(n1430), .Y(n306) );
  NAND2X8TS U500 ( .A(n370), .B(n280), .Y(n403) );
  OAI21X4TS U501 ( .A0(n1915), .A1(n1912), .B0(n1914), .Y(n1909) );
  INVX4TS U502 ( .A(n390), .Y(n493) );
  OAI21X2TS U503 ( .A0(n1834), .A1(n1833), .B0(n136), .Y(n1841) );
  NAND2BX2TS U504 ( .AN(n137), .B(n1828), .Y(n1816) );
  CLKINVX1TS U505 ( .A(n1815), .Y(n137) );
  NAND2X4TS U506 ( .A(n1303), .B(n662), .Y(n363) );
  CLKINVX3TS U507 ( .A(n150), .Y(n149) );
  NOR2BX4TS U508 ( .AN(n1440), .B(n138), .Y(n1445) );
  XOR2X1TS U509 ( .A(n1440), .B(n139), .Y(n1444) );
  NAND2X4TS U510 ( .A(n1303), .B(n787), .Y(n1535) );
  OR2X4TS U511 ( .A(sumOut[59]), .B(n1987), .Y(n275) );
  NAND2X2TS U512 ( .A(n437), .B(n922), .Y(n1493) );
  OAI21X2TS U513 ( .A0(n1296), .A1(n1888), .B0(n1298), .Y(n836) );
  INVX12TS U514 ( .A(n1016), .Y(n991) );
  AOI21X4TS U515 ( .A0(n1843), .A1(n1845), .B0(n919), .Y(n1851) );
  OAI21X4TS U516 ( .A0(n905), .A1(n433), .B0(n446), .Y(n904) );
  INVX16TS U517 ( .A(n192), .Y(n1340) );
  OAI21X2TS U518 ( .A0(n1510), .A1(n2024), .B0(n140), .Y(n1519) );
  AOI21X2TS U519 ( .A0(n1725), .A1(n1729), .B0(n1508), .Y(n140) );
  INVX2TS U520 ( .A(layer2In[2]), .Y(n554) );
  INVX4TS U521 ( .A(n1348), .Y(n1300) );
  OAI2BB1X4TS U522 ( .A0N(n1372), .A1N(n1373), .B0(n142), .Y(n1378) );
  OAI21X4TS U523 ( .A0(n1373), .A1(n1372), .B0(n1370), .Y(n142) );
  XNOR2X4TS U524 ( .A(n264), .B(n147), .Y(n1358) );
  NAND2X8TS U525 ( .A(n1300), .B(n1469), .Y(n147) );
  AND2X8TS U526 ( .A(n1469), .B(n247), .Y(n1465) );
  INVX1TS U527 ( .A(n1728), .Y(n1508) );
  INVX2TS U528 ( .A(n1081), .Y(n1082) );
  INVX6TS U529 ( .A(n1310), .Y(n204) );
  NOR2X6TS U530 ( .A(n178), .B(sumOut[14]), .Y(n1490) );
  XNOR2X4TS U531 ( .A(n960), .B(n966), .Y(n1015) );
  OAI21X4TS U532 ( .A0(n187), .A1(n1259), .B0(sumOut[76]), .Y(n1258) );
  CLKXOR2X4TS U533 ( .A(n1350), .B(n1349), .Y(n1372) );
  CLKINVX3TS U534 ( .A(n145), .Y(n1367) );
  INVX6TS U535 ( .A(n147), .Y(n146) );
  NAND2X2TS U536 ( .A(n1177), .B(weightsIn[58]), .Y(n390) );
  NAND2X4TS U537 ( .A(n184), .B(n1337), .Y(n185) );
  INVX8TS U538 ( .A(n1108), .Y(n1695) );
  NAND2X6TS U539 ( .A(n1313), .B(n1695), .Y(n1323) );
  OAI2BB1X4TS U540 ( .A0N(n1343), .A1N(n301), .B0(n1342), .Y(n1393) );
  NAND2X4TS U541 ( .A(n510), .B(n511), .Y(n319) );
  NOR2X4TS U542 ( .A(n594), .B(n593), .Y(n655) );
  OR2X4TS U543 ( .A(sumOut[29]), .B(n1894), .Y(n270) );
  XOR2X1TS U544 ( .A(n1841), .B(n1840), .Y(genblk1_0__mac_s[9]) );
  INVX2TS U545 ( .A(weightsIn[8]), .Y(n843) );
  XNOR2X4TS U546 ( .A(n150), .B(n893), .Y(n909) );
  NAND2X2TS U547 ( .A(n1469), .B(weightsIn[8]), .Y(n150) );
  INVX6TS U548 ( .A(n554), .Y(n277) );
  OAI21X2TS U549 ( .A0(n1738), .A1(n1744), .B0(n1558), .Y(n759) );
  OR2X8TS U550 ( .A(n472), .B(sumOut[92]), .Y(n2067) );
  XOR2X4TS U551 ( .A(n698), .B(n697), .Y(n700) );
  INVX4TS U552 ( .A(n554), .Y(n566) );
  INVX8TS U553 ( .A(n566), .Y(n358) );
  INVX1TS U554 ( .A(n237), .Y(n630) );
  NAND2X2TS U555 ( .A(n1827), .B(n1828), .Y(n1605) );
  OAI21X4TS U556 ( .A0(n1563), .A1(n1562), .B0(n1561), .Y(n154) );
  NOR2X8TS U557 ( .A(n1478), .B(n1477), .Y(n1563) );
  INVX2TS U558 ( .A(layer2In[0]), .Y(n492) );
  XNOR2X4TS U559 ( .A(n696), .B(n693), .Y(n665) );
  XNOR2X4TS U560 ( .A(n306), .B(n1459), .Y(n1424) );
  OAI21X2TS U561 ( .A0(n1601), .A1(n1833), .B0(n1815), .Y(n1600) );
  XOR2X4TS U562 ( .A(n590), .B(n591), .Y(n569) );
  XNOR2X4TS U563 ( .A(n151), .B(n1201), .Y(n1179) );
  NAND2X8TS U564 ( .A(n1189), .B(n1188), .Y(n151) );
  XOR2X1TS U565 ( .A(n1556), .B(n1555), .Y(genblk1_1__mac_s[7]) );
  XOR2X1TS U566 ( .A(n1488), .B(n1487), .Y(genblk1_1__mac_s[8]) );
  BUFX6TS U567 ( .A(n277), .Y(n1183) );
  INVX6TS U568 ( .A(n492), .Y(n190) );
  NAND2X4TS U569 ( .A(n341), .B(n265), .Y(n340) );
  CLKINVX6TS U570 ( .A(n340), .Y(n1427) );
  NAND2X4TS U571 ( .A(n152), .B(n707), .Y(n681) );
  NAND2X4TS U572 ( .A(n371), .B(n679), .Y(n152) );
  NOR2X4TS U573 ( .A(n594), .B(n1591), .Y(n1612) );
  OR2X4TS U574 ( .A(sumOut[9]), .B(n1838), .Y(n273) );
  XOR2X4TS U575 ( .A(n651), .B(n153), .Y(n600) );
  OAI2BB1X4TS U576 ( .A0N(n590), .A1N(n591), .B0(n589), .Y(n651) );
  NOR2X6TS U577 ( .A(n755), .B(n756), .Y(n945) );
  INVX8TS U578 ( .A(n1016), .Y(n1123) );
  OAI2BB1X4TS U579 ( .A0N(n881), .A1N(n880), .B0(n346), .Y(n935) );
  OAI2BB1X4TS U580 ( .A0N(n1586), .A1N(n1585), .B0(n1584), .Y(n1597) );
  AOI21X4TS U581 ( .A0(n1482), .A1(n1486), .B0(n932), .Y(n933) );
  INVX8TS U582 ( .A(n1177), .Y(n1434) );
  NAND2X4TS U583 ( .A(n425), .B(n1365), .Y(n335) );
  AND2X8TS U584 ( .A(n195), .B(weightsIn[51]), .Y(n1687) );
  NAND2X4TS U585 ( .A(n1177), .B(n1249), .Y(n1209) );
  AOI21X4TS U586 ( .A0(n1566), .A1(n1565), .B0(n154), .Y(n1833) );
  XOR2X4TS U587 ( .A(n1575), .B(n1578), .Y(n344) );
  INVX4TS U588 ( .A(n1603), .Y(n1827) );
  AND2X2TS U589 ( .A(n1827), .B(n1602), .Y(n1599) );
  XOR2X1TS U590 ( .A(n157), .B(n1616), .Y(genblk1_0__mac_s[8]) );
  OAI21X2TS U591 ( .A0(n1605), .A1(n1833), .B0(n1604), .Y(n157) );
  NOR2X8TS U592 ( .A(n1577), .B(n1693), .Y(n1594) );
  INVX4TS U593 ( .A(n195), .Y(n1423) );
  OAI21X4TS U594 ( .A0(n1673), .A1(n1674), .B0(n1671), .Y(n1672) );
  BUFX8TS U595 ( .A(n277), .Y(n1019) );
  OAI21X2TS U596 ( .A0(n1607), .A1(n1608), .B0(sumOut[7]), .Y(n1606) );
  INVX2TS U597 ( .A(n1578), .Y(n1595) );
  XNOR2X4TS U598 ( .A(n160), .B(n1536), .Y(n1541) );
  XOR2X4TS U599 ( .A(n1535), .B(n1539), .Y(n160) );
  OAI21X4TS U600 ( .A0(n1539), .A1(n1538), .B0(n1536), .Y(n1537) );
  XOR2X4TS U601 ( .A(n780), .B(n793), .Y(n812) );
  OAI2BB1X4TS U602 ( .A0N(n799), .A1N(n800), .B0(n779), .Y(n793) );
  OAI21X2TS U603 ( .A0(n1710), .A1(n1982), .B0(n1709), .Y(n1723) );
  AOI21X4TS U604 ( .A0(n1277), .A1(n816), .B0(n815), .Y(n1982) );
  CLKINVX3TS U605 ( .A(n492), .Y(n189) );
  XOR2X4TS U606 ( .A(n801), .B(n161), .Y(n811) );
  XOR2X4TS U607 ( .A(n800), .B(n799), .Y(n161) );
  NAND2X4TS U608 ( .A(n829), .B(n830), .Y(n1707) );
  XOR2X4TS U609 ( .A(n825), .B(n1546), .Y(n829) );
  INVX2TS U610 ( .A(n1542), .Y(n163) );
  OAI2BB1X4TS U611 ( .A0N(n163), .A1N(n162), .B0(n1541), .Y(n294) );
  OAI21X4TS U612 ( .A0(n148), .A1(n1712), .B0(sumOut[57]), .Y(n164) );
  XOR2X4TS U613 ( .A(n1320), .B(n1321), .Y(n179) );
  OAI2BB1X4TS U614 ( .A0N(n1308), .A1N(n1307), .B0(n1306), .Y(n1320) );
  INVX2TS U615 ( .A(n350), .Y(n900) );
  NAND2X4TS U616 ( .A(n1702), .B(n1701), .Y(n1769) );
  OAI2BB1X1TS U617 ( .A0N(n1760), .A1N(n167), .B0(n165), .Y(n1776) );
  XOR2X4TS U618 ( .A(n166), .B(n1760), .Y(n1755) );
  XOR2X4TS U619 ( .A(n1761), .B(n167), .Y(n166) );
  NAND2X4TS U620 ( .A(n1695), .B(n1694), .Y(n167) );
  NOR2X8TS U621 ( .A(n1270), .B(n1269), .Y(n1505) );
  OAI2BB1X4TS U622 ( .A0N(n187), .A1N(n1259), .B0(n1258), .Y(n1270) );
  AOI21X4TS U623 ( .A0(n1792), .A1(n1791), .B0(n1790), .Y(n1793) );
  OAI21X4TS U624 ( .A0(n1770), .A1(n1769), .B0(n1768), .Y(n1792) );
  XOR2X4TS U625 ( .A(n906), .B(sumOut[15]), .Y(n908) );
  NAND2BX4TS U626 ( .AN(n883), .B(n857), .Y(n906) );
  INVX2TS U627 ( .A(n848), .Y(n168) );
  INVX6TS U628 ( .A(n1183), .Y(n745) );
  OAI21X4TS U629 ( .A0(n934), .A1(n1861), .B0(n933), .Y(n943) );
  XOR2X4TS U630 ( .A(n943), .B(n942), .Y(genblk1_1__mac_s[9]) );
  NOR2X6TS U631 ( .A(n814), .B(n813), .Y(n1971) );
  INVX8TS U632 ( .A(n839), .Y(n1633) );
  BUFX6TS U633 ( .A(n298), .Y(n169) );
  BUFX6TS U634 ( .A(n358), .Y(n383) );
  NOR2X8TS U635 ( .A(n465), .B(n241), .Y(n1648) );
  NOR2X4TS U636 ( .A(n222), .B(n171), .Y(n1560) );
  CLKINVX1TS U637 ( .A(n1936), .Y(n1942) );
  OAI21X2TS U638 ( .A0(n552), .A1(n553), .B0(n574), .Y(n286) );
  INVX2TS U639 ( .A(n573), .Y(n552) );
  OAI2BB1X4TS U640 ( .A0N(n577), .A1N(n579), .B0(n559), .Y(n584) );
  OAI2BB1X4TS U641 ( .A0N(n1450), .A1N(n428), .B0(n1435), .Y(n172) );
  BUFX6TS U642 ( .A(n190), .Y(n199) );
  XOR2X4TS U643 ( .A(n1025), .B(n1026), .Y(n173) );
  XOR2X4TS U644 ( .A(n1024), .B(n173), .Y(n1041) );
  NAND2X2TS U645 ( .A(n1025), .B(n1024), .Y(n174) );
  NAND2X2TS U646 ( .A(n170), .B(n1024), .Y(n175) );
  NOR2X8TS U647 ( .A(n1434), .B(n1017), .Y(n1025) );
  OAI21X4TS U648 ( .A0(n1882), .A1(n212), .B0(n353), .Y(n1089) );
  BUFX12TS U649 ( .A(n592), .Y(n877) );
  CLKBUFX2TS U650 ( .A(n1038), .Y(n177) );
  CLKINVX1TS U651 ( .A(n1925), .Y(n1926) );
  XOR2X4TS U652 ( .A(n903), .B(n352), .Y(n178) );
  XNOR2X4TS U653 ( .A(n179), .B(n1315), .Y(n1316) );
  NAND2X4TS U654 ( .A(n1184), .B(n1347), .Y(n1194) );
  OR2X2TS U655 ( .A(n437), .B(n922), .Y(n450) );
  AND2X4TS U656 ( .A(n1177), .B(n1250), .Y(n1190) );
  AND2X8TS U657 ( .A(n199), .B(n968), .Y(n964) );
  INVX8TS U658 ( .A(n839), .Y(n1659) );
  BUFX12TS U659 ( .A(n190), .Y(n839) );
  AND2X4TS U660 ( .A(n839), .B(n1110), .Y(n497) );
  CLKBUFX2TS U661 ( .A(n482), .Y(n180) );
  OAI21X2TS U662 ( .A0(n1466), .A1(n1465), .B0(n1463), .Y(n1464) );
  XNOR2X4TS U663 ( .A(n1645), .B(n1642), .Y(n1624) );
  CLKINVX1TS U664 ( .A(n1642), .Y(n1620) );
  NOR2X4TS U665 ( .A(n1618), .B(n1646), .Y(n1642) );
  INVX4TS U666 ( .A(n200), .Y(n466) );
  NAND2X6TS U667 ( .A(n683), .B(n682), .Y(n716) );
  OAI21X2TS U668 ( .A0(n1917), .A1(n1920), .B0(n1918), .Y(n1901) );
  NAND2X2TS U669 ( .A(sumOut[30]), .B(n1902), .Y(n1920) );
  AND2X2TS U670 ( .A(n991), .B(n853), .Y(n182) );
  AND2X8TS U671 ( .A(n203), .B(n263), .Y(n1344) );
  NAND2X4TS U672 ( .A(n183), .B(n1330), .Y(n186) );
  INVX2TS U673 ( .A(n1337), .Y(n183) );
  INVX4TS U674 ( .A(n1330), .Y(n184) );
  NOR2X6TS U675 ( .A(n1659), .B(n1577), .Y(n1428) );
  XOR2X4TS U676 ( .A(n1255), .B(n1266), .Y(n187) );
  BUFX8TS U677 ( .A(n190), .Y(n1177) );
  AND2X8TS U678 ( .A(n1226), .B(n1225), .Y(n1224) );
  NOR2X4TS U679 ( .A(n1199), .B(sumOut[74]), .Y(n1290) );
  OAI21X2TS U680 ( .A0(n1039), .A1(n1038), .B0(n1037), .Y(n368) );
  OAI21X1TS U681 ( .A0(n2024), .A1(n2023), .B0(n121), .Y(n1273) );
  INVX6TS U682 ( .A(n1347), .Y(n842) );
  AND2X8TS U683 ( .A(n1425), .B(n1019), .Y(n265) );
  INVX4TS U684 ( .A(n592), .Y(n339) );
  AND2X8TS U685 ( .A(n1186), .B(n1185), .Y(n1192) );
  OAI2BB1X2TS U686 ( .A0N(n1681), .A1N(n1680), .B0(n1679), .Y(n1682) );
  BUFX12TS U687 ( .A(n277), .Y(n192) );
  AND2X8TS U688 ( .A(n192), .B(n1351), .Y(n264) );
  AND2X8TS U689 ( .A(n192), .B(n252), .Y(n676) );
  AND2X8TS U690 ( .A(n192), .B(n609), .Y(n610) );
  INVX12TS U691 ( .A(n358), .Y(n195) );
  NOR2X8TS U692 ( .A(n1309), .B(n196), .Y(n1325) );
  BUFX8TS U693 ( .A(n277), .Y(n1347) );
  INVX6TS U694 ( .A(n198), .Y(n1417) );
  INVX6TS U695 ( .A(n1691), .Y(n1635) );
  CLKINVX1TS U696 ( .A(n189), .Y(n188) );
  INVX4TS U697 ( .A(n991), .Y(n594) );
  NOR2X2TS U698 ( .A(n326), .B(n358), .Y(n674) );
  CLKINVX1TS U699 ( .A(n1002), .Y(n1005) );
  CLKINVX1TS U700 ( .A(n398), .Y(n205) );
  INVX2TS U701 ( .A(n205), .Y(n206) );
  CLKAND2X2TS U702 ( .A(n204), .B(n959), .Y(n406) );
  XNOR2X1TS U703 ( .A(n522), .B(n521), .Y(genblk1_9__mac_s[5]) );
  XOR2X4TS U704 ( .A(n673), .B(n672), .Y(n208) );
  INVX2TS U705 ( .A(n1208), .Y(n1213) );
  INVX2TS U706 ( .A(n2009), .Y(n1997) );
  NOR2X4TS U707 ( .A(n2009), .B(n2011), .Y(n722) );
  NOR2X6TS U708 ( .A(n684), .B(sumOut[64]), .Y(n2009) );
  INVX4TS U709 ( .A(n1692), .Y(n1623) );
  INVX4TS U710 ( .A(n305), .Y(n1650) );
  NAND2X4TS U711 ( .A(n478), .B(n477), .Y(n502) );
  OAI2BB1X2TS U712 ( .A0N(n859), .A1N(n858), .B0(n845), .Y(n209) );
  OAI2BB1X2TS U713 ( .A0N(n859), .A1N(n858), .B0(n845), .Y(n872) );
  NAND2X1TS U714 ( .A(n1235), .B(sumOut[74]), .Y(n210) );
  XOR2X1TS U715 ( .A(n1751), .B(n1750), .Y(genblk1_6__mac_s[9]) );
  INVX2TS U716 ( .A(n1880), .Y(n212) );
  NOR2X6TS U717 ( .A(n1647), .B(n1646), .Y(n1688) );
  XOR2X4TS U718 ( .A(n213), .B(n414), .Y(n1199) );
  XOR2X4TS U719 ( .A(n1233), .B(n1231), .Y(n213) );
  OAI21X1TS U720 ( .A0(n1375), .A1(sumOut[35]), .B0(n1316), .Y(n1317) );
  OAI21X4TS U721 ( .A0(n1212), .A1(n1213), .B0(n1210), .Y(n1211) );
  OAI21X2TS U722 ( .A0(n1743), .A1(n1744), .B0(n372), .Y(n1751) );
  NOR2X4TS U723 ( .A(n1658), .B(n358), .Y(n1632) );
  NOR2X4TS U724 ( .A(n923), .B(n922), .Y(n440) );
  OAI2BB1X2TS U725 ( .A0N(n1476), .A1N(n217), .B0(n1474), .Y(n215) );
  NAND2X2TS U726 ( .A(n220), .B(n219), .Y(n221) );
  OR2X2TS U727 ( .A(n1477), .B(n215), .Y(n216) );
  BUFX3TS U728 ( .A(n1490), .Y(n1732) );
  INVX2TS U729 ( .A(n220), .Y(n217) );
  XNOR2X4TS U730 ( .A(n218), .B(n724), .Y(n720) );
  XNOR2X4TS U731 ( .A(n723), .B(sumOut[65]), .Y(n218) );
  NAND2X4TS U732 ( .A(n921), .B(sumOut[14]), .Y(n1491) );
  NAND2X4TS U733 ( .A(n221), .B(n172), .Y(n1474) );
  INVX2TS U734 ( .A(n1476), .Y(n219) );
  INVX2TS U735 ( .A(n1475), .Y(n220) );
  NOR2X4TS U736 ( .A(n1490), .B(n440), .Y(n925) );
  XOR2X4TS U737 ( .A(n1436), .B(n172), .Y(n222) );
  NOR2X4TS U738 ( .A(n383), .B(n843), .Y(n882) );
  OR2X4TS U739 ( .A(n1635), .B(n878), .Y(n863) );
  NOR2X6TS U740 ( .A(n1635), .B(n1205), .Y(n1188) );
  AND2X2TS U741 ( .A(n566), .B(n901), .Y(n899) );
  NAND2X2TS U742 ( .A(n194), .B(n572), .Y(n560) );
  NAND2X2TS U743 ( .A(n198), .B(n1621), .Y(n386) );
  BUFX6TS U744 ( .A(n198), .Y(n1329) );
  INVX1TS U745 ( .A(n1284), .Y(n1285) );
  NAND2X2TS U746 ( .A(n689), .B(n363), .Y(n374) );
  CLKINVX1TS U747 ( .A(n1078), .Y(n1080) );
  XOR2X4TS U748 ( .A(n225), .B(n305), .Y(n1643) );
  XOR2X4TS U749 ( .A(n895), .B(n894), .Y(n897) );
  NOR2X6TS U750 ( .A(n1619), .B(n1646), .Y(n1628) );
  XOR2X1TS U751 ( .A(n336), .B(n2024), .Y(genblk1_7__mac_s[6]) );
  CLKINVX1TS U752 ( .A(n1620), .Y(n223) );
  NOR2X8TS U753 ( .A(n1389), .B(n1390), .Y(n1804) );
  XOR2X4TS U754 ( .A(n351), .B(n1648), .Y(n225) );
  XOR2X4TS U755 ( .A(n230), .B(n514), .Y(n226) );
  OAI21X2TS U756 ( .A0(n1964), .A1(n1967), .B0(n1965), .Y(n1956) );
  NAND2X4TS U757 ( .A(n1161), .B(n1160), .Y(n1528) );
  XNOR2X4TS U758 ( .A(n227), .B(n1755), .Y(n1753) );
  XNOR2X4TS U759 ( .A(n1757), .B(n1758), .Y(n227) );
  XOR2X4TS U760 ( .A(n228), .B(n866), .Y(n873) );
  XOR2X4TS U761 ( .A(n868), .B(n869), .Y(n228) );
  AND2X4TS U762 ( .A(n202), .B(n260), .Y(n498) );
  INVX8TS U763 ( .A(n203), .Y(n1693) );
  OAI21X2TS U764 ( .A0(n1231), .A1(n1233), .B0(n1234), .Y(n1200) );
  CLKINVX1TS U765 ( .A(n2085), .Y(n2086) );
  NOR2X4TS U766 ( .A(n1468), .B(n1577), .Y(n1576) );
  OAI21X1TS U767 ( .A0(n1141), .A1(n1140), .B0(sumOut[97]), .Y(n1139) );
  XOR2X4TS U768 ( .A(n230), .B(n514), .Y(n1152) );
  XNOR2X4TS U769 ( .A(n516), .B(n499), .Y(n230) );
  NOR2X8TS U770 ( .A(n1340), .B(n601), .Y(n611) );
  NOR2X4TS U771 ( .A(n1061), .B(n1060), .Y(n1284) );
  CLKINVX1TS U772 ( .A(n2061), .Y(n2062) );
  XOR2X4TS U773 ( .A(n231), .B(n1260), .Y(n1257) );
  XNOR2X4TS U774 ( .A(n1259), .B(n459), .Y(n231) );
  NAND2X4TS U775 ( .A(n485), .B(n2077), .Y(n1158) );
  NAND2X4TS U776 ( .A(n1163), .B(n1162), .Y(n1530) );
  XNOR2X4TS U777 ( .A(n488), .B(n510), .Y(n495) );
  BUFX6TS U778 ( .A(layer2In[3]), .Y(n592) );
  INVX2TS U779 ( .A(n1357), .Y(n232) );
  CLKINVX3TS U780 ( .A(n232), .Y(n233) );
  OAI2BB1X4TS U781 ( .A0N(n733), .A1N(n732), .B0(n731), .Y(n744) );
  OAI21X2TS U782 ( .A0(n406), .A1(n966), .B0(n964), .Y(n965) );
  XOR2X4TS U783 ( .A(n782), .B(n781), .Y(n234) );
  OAI2BB1X2TS U784 ( .A0N(n581), .A1N(n457), .B0(n637), .Y(n582) );
  NAND2X2TS U785 ( .A(n1019), .B(n1018), .Y(n235) );
  XOR2X4TS U786 ( .A(n234), .B(n783), .Y(n236) );
  NOR2X4TS U787 ( .A(n1633), .B(n1534), .Y(n783) );
  OAI21X1TS U788 ( .A0(sumOut[15]), .A1(n906), .B0(n447), .Y(n861) );
  NOR2X4TS U789 ( .A(n920), .B(sumOut[13]), .Y(n1848) );
  XOR2X1TS U790 ( .A(n624), .B(n623), .Y(n237) );
  OAI21X2TS U791 ( .A0(n1573), .A1(n1572), .B0(n1570), .Y(n1571) );
  NAND2X2TS U792 ( .A(n645), .B(n644), .Y(n1298) );
  NAND2X2TS U793 ( .A(n395), .B(n1384), .Y(n1927) );
  XOR2X4TS U794 ( .A(n238), .B(n1685), .Y(n1679) );
  XOR2X4TS U795 ( .A(n1688), .B(n1687), .Y(n238) );
  NAND2X4TS U796 ( .A(n1691), .B(n1250), .Y(n1208) );
  INVX2TS U797 ( .A(n200), .Y(n239) );
  NOR2X4TS U798 ( .A(n1434), .B(n1421), .Y(n1447) );
  NOR2X4TS U799 ( .A(n1434), .B(n1591), .Y(n1463) );
  NOR2X2TS U800 ( .A(n1434), .B(n364), .Y(n1656) );
  NOR2X4TS U801 ( .A(n678), .B(n326), .Y(n701) );
  NOR2X2TS U802 ( .A(n244), .B(n1658), .Y(n2042) );
  AND2X4TS U803 ( .A(n668), .B(n969), .Y(n677) );
  CLKINVX6TS U804 ( .A(n1690), .Y(n240) );
  CLKINVX1TS U805 ( .A(n240), .Y(n242) );
  CLKINVX1TS U806 ( .A(n240), .Y(n243) );
  INVX6TS U807 ( .A(n969), .Y(n1619) );
  CLKINVX1TS U808 ( .A(n194), .Y(n245) );
  NOR2X2TS U809 ( .A(n1715), .B(n838), .Y(n881) );
  OR2X4TS U810 ( .A(n245), .B(n1779), .Y(n1798) );
  NAND2X4TS U811 ( .A(n1303), .B(n1252), .Y(n332) );
  NAND2X4TS U812 ( .A(n1691), .B(n766), .Y(n782) );
  NAND2X2TS U813 ( .A(n204), .B(n255), .Y(n299) );
  NAND2X4TS U814 ( .A(n204), .B(n1426), .Y(n304) );
  CLKINVX1TS U815 ( .A(n887), .Y(n246) );
  INVX4TS U816 ( .A(n1577), .Y(n247) );
  INVX2TS U817 ( .A(n656), .Y(n248) );
  INVX2TS U818 ( .A(weightsIn[19]), .Y(n249) );
  CLKINVX3TS U819 ( .A(n249), .Y(n250) );
  CLKINVX1TS U820 ( .A(n249), .Y(n251) );
  INVX2TS U821 ( .A(n703), .Y(n252) );
  CLKINVX3TS U822 ( .A(weightsIn[44]), .Y(n253) );
  INVX2TS U823 ( .A(n253), .Y(n254) );
  CLKINVX1TS U824 ( .A(n253), .Y(n255) );
  INVX2TS U825 ( .A(n256), .Y(n257) );
  CLKINVX1TS U826 ( .A(n256), .Y(n258) );
  INVX2TS U827 ( .A(weightsIn[21]), .Y(n261) );
  INVX2TS U828 ( .A(n261), .Y(n262) );
  CLKINVX1TS U829 ( .A(n261), .Y(n263) );
  OAI21X1TS U830 ( .A0(n1410), .A1(n1411), .B0(sumOut[38]), .Y(n322) );
  OAI2BB1X2TS U831 ( .A0N(n894), .A1N(n895), .B0(n891), .Y(n905) );
  XOR2X1TS U832 ( .A(n1411), .B(sumOut[38]), .Y(n323) );
  XOR2X1TS U833 ( .A(n1410), .B(n323), .Y(n1399) );
  OAI21X1TS U834 ( .A0(n1874), .A1(n1877), .B0(n1875), .Y(n1866) );
  NAND2X1TS U835 ( .A(sumOut[80]), .B(n2042), .Y(n2056) );
  NAND2X1TS U836 ( .A(n1919), .B(n1918), .Y(n1921) );
  AND2X4TS U837 ( .A(n1313), .B(n200), .Y(n266) );
  INVX2TS U838 ( .A(n663), .Y(n281) );
  BUFX8TS U839 ( .A(n465), .Y(n1214) );
  AND2X4TS U840 ( .A(n969), .B(n572), .Y(n267) );
  OR2X2TS U841 ( .A(sumOut[89]), .B(n1800), .Y(n268) );
  OR2X1TS U842 ( .A(sumOut[69]), .B(n1748), .Y(n269) );
  XOR2X4TS U843 ( .A(n859), .B(n858), .Y(n444) );
  OR2X1TS U844 ( .A(sumOut[99]), .B(n1173), .Y(n271) );
  OR2X2TS U845 ( .A(sumOut[39]), .B(n1413), .Y(n272) );
  NAND2X4TS U846 ( .A(n718), .B(sumOut[64]), .Y(n398) );
  INVX1TS U847 ( .A(n1276), .Y(n411) );
  CLKINVX2TS U848 ( .A(n1817), .Y(n1819) );
  INVX1TS U849 ( .A(n1943), .Y(n1944) );
  NAND2X2TS U850 ( .A(n1721), .B(n1720), .Y(n1977) );
  CLKINVX2TS U851 ( .A(n2080), .Y(n2082) );
  XOR2X1TS U852 ( .A(n1170), .B(n1151), .Y(n1164) );
  CLKINVX2TS U853 ( .A(n1336), .Y(n1333) );
  INVX2TS U854 ( .A(n1783), .Y(n1781) );
  CLKINVX2TS U855 ( .A(n1959), .Y(n1961) );
  OAI2BB1X2TS U856 ( .A0N(n1149), .A1N(n1148), .B0(n1147), .Y(n1170) );
  INVX1TS U857 ( .A(n2033), .Y(n2035) );
  CLKINVX1TS U858 ( .A(n1948), .Y(n1950) );
  INVX1TS U859 ( .A(n1917), .Y(n1919) );
  CLKINVX2TS U860 ( .A(n798), .Y(n795) );
  INVX1TS U861 ( .A(n2004), .Y(n2006) );
  INVX2TS U862 ( .A(n403), .Y(n366) );
  OAI21X2TS U863 ( .A0(n1718), .A1(n1719), .B0(n1716), .Y(n1717) );
  INVX1TS U864 ( .A(n2053), .Y(n2055) );
  OAI21X2TS U865 ( .A0(n1446), .A1(n1447), .B0(n1445), .Y(n377) );
  INVX2TS U866 ( .A(n1853), .Y(n1855) );
  NAND2X4TS U867 ( .A(n688), .B(n424), .Y(n292) );
  INVX3TS U868 ( .A(n706), .Y(n371) );
  NOR2X4TS U869 ( .A(n332), .B(n329), .Y(n331) );
  INVX1TS U870 ( .A(n880), .Y(n348) );
  INVX3TS U871 ( .A(n342), .Y(n341) );
  XOR2X1TS U872 ( .A(sumOut[98]), .B(n1171), .Y(n1151) );
  INVX3TS U873 ( .A(n424), .Y(n689) );
  INVX2TS U874 ( .A(n456), .Y(n449) );
  BUFX3TS U875 ( .A(weightsIn[33]), .Y(n766) );
  BUFX4TS U876 ( .A(weightsIn[13]), .Y(n282) );
  INVX1TS U877 ( .A(n1765), .Y(n1766) );
  AND2X2TS U878 ( .A(n271), .B(n1174), .Y(n1175) );
  XOR2X1TS U879 ( .A(n1278), .B(n1970), .Y(genblk1_5__mac_s[4]) );
  INVX1TS U880 ( .A(n1524), .Y(n1166) );
  INVX1TS U881 ( .A(n1518), .Y(n379) );
  INVX2TS U882 ( .A(n1831), .Y(n1604) );
  CLKINVX2TS U883 ( .A(n1886), .Y(n648) );
  NAND2BX2TS U884 ( .AN(n2023), .B(n121), .Y(n336) );
  INVX2TS U885 ( .A(n1529), .Y(n1531) );
  NOR2X2TS U886 ( .A(n832), .B(n1296), .Y(n1883) );
  INVX1TS U887 ( .A(n1094), .Y(n1066) );
  XOR2X1TS U888 ( .A(n2084), .B(n2083), .Y(genblk1_9__mac_s[1]) );
  NOR2X4TS U889 ( .A(n646), .B(n647), .Y(n832) );
  OAI2BB1X1TS U890 ( .A0N(n1171), .A1N(n1170), .B0(n1169), .Y(n1172) );
  NAND2X1TS U891 ( .A(n2082), .B(n2081), .Y(n2084) );
  XOR2X1TS U892 ( .A(n2037), .B(n2036), .Y(genblk1_7__mac_s[1]) );
  NAND2X4TS U893 ( .A(n1248), .B(n1247), .Y(n1259) );
  NAND2X2TS U894 ( .A(sumOut[92]), .B(n472), .Y(n2066) );
  NAND2X4TS U895 ( .A(n695), .B(n285), .Y(n723) );
  OAI2BB1X2TS U896 ( .A0N(n1411), .A1N(n1410), .B0(n322), .Y(n1412) );
  XOR2X1TS U897 ( .A(n1952), .B(n1951), .Y(genblk1_4__mac_s[1]) );
  AOI21X2TS U898 ( .A0(n2039), .A1(n2041), .B0(n1662), .Y(n2051) );
  INVX1TS U899 ( .A(n1930), .Y(n1054) );
  XOR2X1TS U900 ( .A(n1878), .B(n1877), .Y(genblk1_2__mac_s[1]) );
  INVX1TS U901 ( .A(n1809), .Y(n1449) );
  XOR2X1TS U902 ( .A(n2057), .B(n2056), .Y(genblk1_8__mac_s[1]) );
  NAND2X1TS U903 ( .A(n1950), .B(n1949), .Y(n1952) );
  XOR2X1TS U904 ( .A(n1968), .B(n1967), .Y(genblk1_5__mac_s[1]) );
  XOR2X1TS U905 ( .A(n2008), .B(n2007), .Y(genblk1_6__mac_s[1]) );
  NAND2XLTS U906 ( .A(n2055), .B(n2054), .Y(n2057) );
  NAND2XLTS U907 ( .A(n1966), .B(n1965), .Y(n1968) );
  OAI2BB1X1TS U908 ( .A0N(n1892), .A1N(n1891), .B0(n1890), .Y(n1893) );
  NAND2X2TS U909 ( .A(sumOut[72]), .B(n1228), .Y(n2016) );
  NAND2X2TS U910 ( .A(sumOut[12]), .B(n918), .Y(n1842) );
  NAND2XLTS U911 ( .A(n1824), .B(n1823), .Y(n1826) );
  NAND2XLTS U912 ( .A(n2006), .B(n2005), .Y(n2008) );
  NAND2X2TS U913 ( .A(sumOut[32]), .B(n1360), .Y(n1898) );
  NAND2XLTS U914 ( .A(n1876), .B(n1875), .Y(n1878) );
  XOR2X1TS U915 ( .A(n1857), .B(n1856), .Y(genblk1_1__mac_s[1]) );
  INVX3TS U916 ( .A(n1231), .Y(n1232) );
  INVX1TS U917 ( .A(n634), .Y(n631) );
  NAND2X4TS U918 ( .A(n292), .B(n374), .Y(n664) );
  NAND2X1TS U919 ( .A(n1855), .B(n1854), .Y(n1857) );
  INVX1TS U920 ( .A(n1874), .Y(n1876) );
  INVX1TS U921 ( .A(n1822), .Y(n1824) );
  CLKBUFX2TS U922 ( .A(n106), .Y(n550) );
  AND2X2TS U923 ( .A(n1903), .B(n1920), .Y(genblk1_3__mac_s[0]) );
  XOR2X1TS U924 ( .A(n1891), .B(n657), .Y(n658) );
  CLKBUFX2TS U925 ( .A(n22), .Y(n551) );
  AND2X2TS U926 ( .A(n1814), .B(n1825), .Y(genblk1_0__mac_s[0]) );
  AND2X2TS U927 ( .A(n1935), .B(n1951), .Y(genblk1_4__mac_s[0]) );
  OAI21X1TS U928 ( .A0(n1891), .A1(n1892), .B0(sumOut[28]), .Y(n1890) );
  CLKBUFX2TS U929 ( .A(n540), .Y(n541) );
  CLKBUFX2TS U930 ( .A(n543), .Y(n544) );
  CLKBUFX2TS U931 ( .A(n528), .Y(n529) );
  CLKBUFX2TS U932 ( .A(n526), .Y(n527) );
  CLKBUFX2TS U933 ( .A(n70), .Y(n547) );
  CLKBUFX2TS U934 ( .A(n548), .Y(n549) );
  CLKBUFX2TS U935 ( .A(n45), .Y(n530) );
  NAND2X2TS U936 ( .A(sumOut[40]), .B(n1934), .Y(n1951) );
  INVX2TS U937 ( .A(n1663), .Y(n1664) );
  CLKBUFX2TS U938 ( .A(n531), .Y(n532) );
  CLKBUFX2TS U939 ( .A(n10), .Y(n542) );
  AND2X2TS U940 ( .A(n2021), .B(n2036), .Y(genblk1_7__mac_s[0]) );
  INVX1TS U941 ( .A(n881), .Y(n347) );
  ADDFHX2TS U942 ( .A(n655), .B(n654), .CI(n653), .CO(n1891), .S(n652) );
  INVX2TS U943 ( .A(n715), .Y(n278) );
  INVX3TS U944 ( .A(n1315), .Y(n1318) );
  CLKBUFX2TS U945 ( .A(n537), .Y(n538) );
  AND2X2TS U946 ( .A(n1958), .B(n1967), .Y(genblk1_5__mac_s[0]) );
  AND2X4TS U947 ( .A(n1049), .B(n1048), .Y(n1046) );
  CLKBUFX2TS U948 ( .A(n105), .Y(n536) );
  CLKBUFX2TS U949 ( .A(n94), .Y(n545) );
  CLKBUFX2TS U950 ( .A(n118), .Y(n546) );
  CLKBUFX2TS U951 ( .A(n523), .Y(n524) );
  OR2X2TS U952 ( .A(sumOut[70]), .B(n2020), .Y(n2021) );
  AND2X2TS U953 ( .A(n1995), .B(n2007), .Y(genblk1_6__mac_s[0]) );
  OR2X2TS U954 ( .A(n1715), .B(n951), .Y(n1746) );
  AND2X2TS U955 ( .A(n2071), .B(n2083), .Y(genblk1_9__mac_s[0]) );
  INVX1TS U956 ( .A(n591), .Y(n588) );
  AND2X2TS U957 ( .A(n1868), .B(n1877), .Y(genblk1_2__mac_s[0]) );
  CLKBUFX2TS U958 ( .A(n81), .Y(n525) );
  NAND2X4TS U959 ( .A(n1123), .B(n901), .Y(n888) );
  INVX1TS U960 ( .A(n1634), .Y(n387) );
  INVX1TS U961 ( .A(n1321), .Y(n314) );
  INVX1TS U962 ( .A(n1684), .Y(n1680) );
  INVX1TS U963 ( .A(n894), .Y(n890) );
  CLKBUFX2TS U964 ( .A(n533), .Y(n534) );
  INVX2TS U965 ( .A(sumOut[35]), .Y(n1374) );
  INVX2TS U966 ( .A(sumOut[62]), .Y(n710) );
  INVX2TS U967 ( .A(sumOut[47]), .Y(n993) );
  INVX1TS U968 ( .A(sumOut[96]), .Y(n439) );
  INVX2TS U969 ( .A(n1499), .Y(n1252) );
  CLKINVX2TS U970 ( .A(n1779), .Y(n1694) );
  CLKINVX2TS U971 ( .A(n951), .Y(n735) );
  INVX2TS U972 ( .A(n1180), .Y(n1184) );
  INVX4TS U973 ( .A(n766), .Y(n823) );
  INVX2TS U974 ( .A(n1029), .Y(n280) );
  INVX1TS U975 ( .A(weightsIn[31]), .Y(n776) );
  BUFX3TS U976 ( .A(weightsIn[31]), .Y(n767) );
  INVX2TS U977 ( .A(weightsIn[6]), .Y(n887) );
  AOI21X4TS U978 ( .A0(n1238), .A1(n1289), .B0(n283), .Y(n2024) );
  OAI21X4TS U979 ( .A0(n1291), .A1(n1292), .B0(n1293), .Y(n283) );
  NAND2X4TS U980 ( .A(n1691), .B(n281), .Y(n730) );
  AND2X8TS U981 ( .A(n455), .B(n461), .Y(n772) );
  OAI21X4TS U982 ( .A0(n1529), .A1(n1528), .B0(n1530), .Y(n1521) );
  OAI2BB1X4TS U983 ( .A0N(n743), .A1N(n744), .B0(n742), .Y(n949) );
  AND2X4TS U984 ( .A(n281), .B(n198), .Y(n750) );
  OAI21X4TS U985 ( .A0(n945), .A1(n1558), .B0(n944), .Y(n1742) );
  NOR2X8TS U986 ( .A(n1693), .B(n1442), .Y(n1429) );
  OAI2BB1X2TS U987 ( .A0N(n553), .A1N(n552), .B0(n286), .Y(n579) );
  AND2X8TS U988 ( .A(n774), .B(n384), .Y(n791) );
  XOR2X4TS U989 ( .A(n827), .B(n408), .Y(n814) );
  OAI21X2TS U990 ( .A0(n1982), .A1(n1705), .B0(n130), .Y(n1551) );
  INVX4TS U991 ( .A(n199), .Y(n898) );
  OAI21X4TS U992 ( .A0(n804), .A1(n802), .B0(n803), .Y(n778) );
  OAI21X4TS U993 ( .A0(n394), .A1(n1547), .B0(sumOut[56]), .Y(n1545) );
  XNOR2X4TS U994 ( .A(n289), .B(n1541), .Y(n394) );
  XNOR2X4TS U995 ( .A(n1542), .B(n1543), .Y(n289) );
  NAND2X4TS U996 ( .A(n291), .B(n290), .Y(n826) );
  CLKINVX1TS U997 ( .A(n791), .Y(n290) );
  NAND2X4TS U998 ( .A(n789), .B(n236), .Y(n291) );
  INVX2TS U999 ( .A(n729), .Y(n690) );
  XOR2X4TS U1000 ( .A(n293), .B(n1541), .Y(n1546) );
  XOR2X4TS U1001 ( .A(n1542), .B(n1543), .Y(n293) );
  AND2X8TS U1002 ( .A(n202), .B(n837), .Y(n460) );
  XNOR2X4TS U1003 ( .A(n732), .B(n730), .Y(n362) );
  NOR2X8TS U1004 ( .A(n383), .B(n1181), .Y(n1189) );
  XOR2X4TS U1005 ( .A(n295), .B(n911), .Y(n920) );
  NOR2X4TS U1006 ( .A(n1128), .B(n1129), .Y(n1144) );
  NAND2X4TS U1007 ( .A(n1257), .B(n1256), .Y(n2022) );
  OAI2BB1X4TS U1008 ( .A0N(n169), .A1N(n1254), .B0(n296), .Y(n1266) );
  OAI21X4TS U1009 ( .A0(n1254), .A1(n169), .B0(n1253), .Y(n296) );
  XOR2X4TS U1010 ( .A(n297), .B(n1254), .Y(n1242) );
  XOR2X4TS U1011 ( .A(n1253), .B(n298), .Y(n297) );
  XOR2X4TS U1012 ( .A(n300), .B(n330), .Y(n1264) );
  XOR2X4TS U1013 ( .A(n329), .B(n356), .Y(n300) );
  OR2X4TS U1014 ( .A(n134), .B(n656), .Y(n654) );
  OAI2BB1X2TS U1015 ( .A0N(n916), .A1N(n915), .B0(n302), .Y(n911) );
  XNOR2X4TS U1016 ( .A(n303), .B(n914), .Y(n918) );
  XNOR2X4TS U1017 ( .A(n915), .B(n916), .Y(n303) );
  NAND2X4TS U1018 ( .A(n1461), .B(n306), .Y(n1569) );
  INVX2TS U1019 ( .A(n1884), .Y(n1885) );
  XOR2X4TS U1020 ( .A(n1465), .B(n1466), .Y(n1419) );
  OAI21X2TS U1021 ( .A0(n1629), .A1(n1639), .B0(n458), .Y(n1638) );
  NAND2X4TS U1022 ( .A(n1623), .B(n198), .Y(n305) );
  XOR2X4TS U1023 ( .A(n1430), .B(n307), .Y(n1450) );
  ADDFHX4TS U1024 ( .A(n615), .B(n614), .CI(n613), .CO(n618), .S(n607) );
  XNOR2X4TS U1025 ( .A(n309), .B(n1098), .Y(n1115) );
  XOR2X4TS U1026 ( .A(n1099), .B(n1102), .Y(n309) );
  OAI21X2TS U1027 ( .A0(n1889), .A1(n1888), .B0(n312), .Y(n1897) );
  AOI21X4TS U1028 ( .A0(n1886), .A1(n1887), .B0(n1885), .Y(n312) );
  OAI2BB1X4TS U1029 ( .A0N(n314), .A1N(n313), .B0(n1318), .Y(n1319) );
  XOR2X4TS U1030 ( .A(n317), .B(n474), .Y(n472) );
  NAND2X4TS U1031 ( .A(n319), .B(n318), .Y(n1118) );
  OAI21X4TS U1032 ( .A0(n1906), .A1(n1804), .B0(n1806), .Y(n1407) );
  NAND2X4TS U1033 ( .A(n321), .B(n320), .Y(n1397) );
  NOR2X4TS U1034 ( .A(n1230), .B(sumOut[73]), .Y(n2028) );
  INVX2TS U1035 ( .A(n1181), .Y(n1182) );
  OAI2BB1X4TS U1036 ( .A0N(n1212), .A1N(n1213), .B0(n1211), .Y(n1245) );
  NOR2X8TS U1037 ( .A(n1693), .B(n1181), .Y(n1212) );
  AND2X2TS U1038 ( .A(n1406), .B(n1404), .Y(n1401) );
  OAI21X4TS U1039 ( .A0(n1298), .A1(n832), .B0(n833), .Y(n1886) );
  NAND2X2TS U1040 ( .A(n920), .B(sumOut[13]), .Y(n1850) );
  XOR2X4TS U1041 ( .A(n1569), .B(sumOut[5]), .Y(n1472) );
  XOR2X4TS U1042 ( .A(n1364), .B(n1363), .Y(n1366) );
  OAI2BB1X4TS U1043 ( .A0N(n1335), .A1N(n1336), .B0(n1334), .Y(n1389) );
  INVX4TS U1044 ( .A(n198), .Y(n1207) );
  XOR2X4TS U1045 ( .A(n666), .B(n278), .Y(n717) );
  INVX2TS U1046 ( .A(n257), .Y(n326) );
  INVX2TS U1047 ( .A(n332), .Y(n330) );
  OAI2BB2X4TS U1048 ( .B0(n331), .B1(n135), .A0N(n329), .A1N(n332), .Y(n1500)
         );
  OAI21X1TS U1049 ( .A0(n1502), .A1(n1503), .B0(n1500), .Y(n1501) );
  INVX2TS U1050 ( .A(n334), .Y(n553) );
  XOR2X4TS U1051 ( .A(n573), .B(n334), .Y(n575) );
  XOR2X4TS U1052 ( .A(n803), .B(n802), .Y(n805) );
  OAI2BB1X4TS U1053 ( .A0N(n747), .A1N(n357), .B0(n746), .Y(n748) );
  XOR2X4TS U1054 ( .A(n375), .B(n337), .Y(n1304) );
  NAND2X4TS U1055 ( .A(n1300), .B(n193), .Y(n337) );
  NOR2X4TS U1056 ( .A(n1598), .B(n1597), .Y(n1603) );
  ADDFHX4TS U1057 ( .A(n498), .B(n497), .CI(n496), .CO(n517), .S(n500) );
  INVX2TS U1058 ( .A(n517), .Y(n499) );
  NOR2X4TS U1059 ( .A(n830), .B(n829), .Y(n1705) );
  XOR2X4TS U1060 ( .A(n1629), .B(n1639), .Y(n1630) );
  NOR2X8TS U1061 ( .A(n1658), .B(n1625), .Y(n1639) );
  NOR2X2TS U1062 ( .A(sumOut[41]), .B(n1052), .Y(n1948) );
  NAND2X2TS U1063 ( .A(n419), .B(n1279), .Y(n1283) );
  XOR2X1TS U1064 ( .A(n1897), .B(n1896), .Y(genblk1_2__mac_s[9]) );
  NOR2X4TS U1065 ( .A(n812), .B(sumOut[54]), .Y(n1274) );
  AND2X2TS U1066 ( .A(n1095), .B(n1094), .Y(n1096) );
  XOR2X1TS U1067 ( .A(n605), .B(n606), .Y(n603) );
  OAI21X4TS U1068 ( .A0(n620), .A1(n619), .B0(n618), .Y(n355) );
  XNOR2X4TS U1069 ( .A(n265), .B(n342), .Y(n1446) );
  INVX2TS U1070 ( .A(n1653), .Y(n343) );
  OAI2BB1X4TS U1071 ( .A0N(n1634), .A1N(n343), .B0(n385), .Y(n1666) );
  OAI2BB1X4TS U1072 ( .A0N(n460), .A1N(n854), .B0(n840), .Y(n859) );
  XOR2X4TS U1073 ( .A(n344), .B(n1576), .Y(n1570) );
  NOR2X8TS U1074 ( .A(n345), .B(n1676), .Y(n2061) );
  XOR2X4TS U1075 ( .A(n1652), .B(n1698), .Y(n1676) );
  OAI2BB1X4TS U1076 ( .A0N(n1674), .A1N(n1673), .B0(n1641), .Y(n345) );
  NOR2X4TS U1077 ( .A(n2023), .B(n1505), .Y(n1724) );
  INVX2TS U1078 ( .A(n1724), .Y(n1727) );
  AND2X4TS U1079 ( .A(n1695), .B(n246), .Y(n912) );
  OAI2BB1X2TS U1080 ( .A0N(n348), .A1N(n347), .B0(n879), .Y(n346) );
  XOR2X4TS U1081 ( .A(n876), .B(sumOut[17]), .Y(n870) );
  XNOR2X4TS U1082 ( .A(n349), .B(n879), .Y(n876) );
  XNOR2X4TS U1083 ( .A(n881), .B(n880), .Y(n349) );
  OAI21X2TS U1084 ( .A0(n585), .A1(n584), .B0(sumOut[26]), .Y(n583) );
  XNOR2X4TS U1085 ( .A(n350), .B(n899), .Y(n915) );
  INVX2TS U1086 ( .A(n1802), .Y(n378) );
  INVX4TS U1087 ( .A(n1770), .Y(n1787) );
  OAI21X4TS U1088 ( .A0(n1343), .A1(n301), .B0(n1341), .Y(n1342) );
  OAI21X4TS U1089 ( .A0(n799), .A1(n800), .B0(n801), .Y(n779) );
  OAI2BB1X4TS U1090 ( .A0N(n802), .A1N(n804), .B0(n778), .Y(n801) );
  NOR2X4TS U1091 ( .A(n1256), .B(n1257), .Y(n2023) );
  AND2X2TS U1092 ( .A(n1887), .B(n1884), .Y(n660) );
  XOR2X4TS U1093 ( .A(n903), .B(n352), .Y(n921) );
  OAI2BB1X4TS U1094 ( .A0N(n910), .A1N(n909), .B0(n902), .Y(n352) );
  BUFX3TS U1095 ( .A(n1084), .Y(n353) );
  CLKINVX1TS U1096 ( .A(n483), .Y(n2078) );
  NAND2BX4TS U1097 ( .AN(n473), .B(n354), .Y(n483) );
  XNOR2X2TS U1098 ( .A(n1089), .B(n1088), .Y(genblk1_2__mac_s[5]) );
  OAI2BB1X4TS U1099 ( .A0N(n620), .A1N(n619), .B0(n355), .Y(n629) );
  NOR2X4TS U1100 ( .A(n1290), .B(n1292), .Y(n1238) );
  NOR2X6TS U1101 ( .A(n1237), .B(n1236), .Y(n1292) );
  XOR2X1TS U1102 ( .A(n1273), .B(n1272), .Y(genblk1_7__mac_s[7]) );
  XOR2X4TS U1103 ( .A(n1208), .B(n1209), .Y(n1178) );
  CLKBUFX2TS U1104 ( .A(n693), .Y(n359) );
  XOR2X4TS U1105 ( .A(n360), .B(n233), .Y(n1360) );
  OAI2BB1X2TS U1106 ( .A0N(n1398), .A1N(n1397), .B0(n1396), .Y(n1400) );
  XNOR2X4TS U1107 ( .A(n362), .B(n733), .Y(n726) );
  OAI21X4TS U1108 ( .A0(n2061), .A1(n2045), .B0(n2063), .Y(n1677) );
  CLKINVX3TS U1109 ( .A(n797), .Y(n794) );
  INVX2TS U1110 ( .A(n794), .Y(n427) );
  XOR2X4TS U1111 ( .A(n862), .B(n865), .Y(n404) );
  OAI21X2TS U1112 ( .A0(n980), .A1(n979), .B0(n985), .Y(n978) );
  XOR2X4TS U1113 ( .A(n1314), .B(n1323), .Y(n1315) );
  NAND2X4TS U1114 ( .A(n359), .B(n694), .Y(n695) );
  NOR2X4TS U1115 ( .A(n2085), .B(n1529), .Y(n1520) );
  NOR2X8TS U1116 ( .A(n1162), .B(n1163), .Y(n1529) );
  NOR2X4TS U1117 ( .A(n1635), .B(n1180), .Y(n1225) );
  AND2X8TS U1118 ( .A(n1628), .B(n365), .Y(n1645) );
  XOR2X4TS U1119 ( .A(n365), .B(n1628), .Y(n1663) );
  NOR2X8TS U1120 ( .A(n1618), .B(n364), .Y(n365) );
  AOI21X4TS U1121 ( .A0(n1059), .A1(n1936), .B0(n367), .Y(n1287) );
  OAI21X4TS U1122 ( .A0(n1280), .A1(n1937), .B0(n1281), .Y(n367) );
  OAI21X4TS U1123 ( .A0(n1307), .A1(n1308), .B0(n266), .Y(n1306) );
  OAI2BB1X4TS U1124 ( .A0N(n1039), .A1N(n177), .B0(n368), .Y(n1057) );
  OAI21X4TS U1125 ( .A0(n1795), .A1(n1794), .B0(n1793), .Y(n1803) );
  XOR2X4TS U1126 ( .A(n1803), .B(n378), .Y(genblk1_8__mac_s[9]) );
  NOR2X4TS U1127 ( .A(n1017), .B(n1326), .Y(n979) );
  XOR2X4TS U1128 ( .A(n1590), .B(n156), .Y(n1580) );
  OAI2BB1X4TS U1129 ( .A0N(n1576), .A1N(n1575), .B0(n1574), .Y(n1590) );
  NAND2X4TS U1130 ( .A(n258), .B(n204), .Y(n424) );
  XNOR2X4TS U1131 ( .A(n1014), .B(n403), .Y(n402) );
  CLKINVX1TS U1132 ( .A(n666), .Y(n423) );
  OAI2BB1X4TS U1133 ( .A0N(n278), .A1N(n666), .B0(n716), .Y(n685) );
  NAND2X4TS U1134 ( .A(n740), .B(n739), .Y(n1558) );
  AOI21X4TS U1135 ( .A0(n1742), .A1(n1741), .B0(n1740), .Y(n372) );
  NOR2X8TS U1136 ( .A(n1468), .B(n734), .Y(n732) );
  AND2X2TS U1137 ( .A(n1554), .B(n1553), .Y(n1555) );
  NAND2X2TS U1138 ( .A(n793), .B(n373), .Y(n796) );
  NAND2X2TS U1139 ( .A(n794), .B(n795), .Y(n373) );
  OAI21X2TS U1140 ( .A0(n2085), .A1(n2087), .B0(n1528), .Y(n1533) );
  XOR2X4TS U1141 ( .A(n481), .B(n207), .Y(n484) );
  XOR2X4TS U1142 ( .A(n635), .B(sumOut[25]), .Y(n636) );
  NAND2BX4TS U1143 ( .AN(n622), .B(n576), .Y(n635) );
  XOR2X4TS U1144 ( .A(n376), .B(n1445), .Y(n1448) );
  XOR2X4TS U1145 ( .A(n1446), .B(n1447), .Y(n376) );
  OAI21X4TS U1146 ( .A0(n1451), .A1(n1450), .B0(n1452), .Y(n1435) );
  OAI2BB1X4TS U1147 ( .A0N(n1001), .A1N(n1000), .B0(n999), .Y(n1062) );
  INVX2TS U1148 ( .A(n1285), .Y(n410) );
  XOR2X1TS U1149 ( .A(n1519), .B(n379), .Y(genblk1_7__mac_s[9]) );
  XOR2X4TS U1150 ( .A(n380), .B(n1341), .Y(n1337) );
  XNOR2X4TS U1151 ( .A(n1323), .B(n1344), .Y(n380) );
  OAI2BB1X4TS U1152 ( .A0N(n1324), .A1N(n1325), .B0(n382), .Y(n1339) );
  XOR2X4TS U1153 ( .A(n774), .B(n384), .Y(n799) );
  NOR2X4TS U1154 ( .A(n196), .B(n776), .Y(n384) );
  OAI2BB1X4TS U1155 ( .A0N(n387), .A1N(n1653), .B0(n1654), .Y(n385) );
  XOR2X4TS U1156 ( .A(n386), .B(n1632), .Y(n1653) );
  NOR2X8TS U1157 ( .A(n466), .B(n734), .Y(n670) );
  NOR2X1TS U1158 ( .A(n466), .B(n703), .Y(n1994) );
  AOI2BB2X4TS U1159 ( .B0(n389), .B1(n493), .A0N(n338), .A1N(n388), .Y(n1099)
         );
  OAI2BB1X4TS U1160 ( .A0N(n818), .A1N(n393), .B0(n391), .Y(n1547) );
  OAI21X4TS U1161 ( .A0(n818), .A1(n393), .B0(n817), .Y(n391) );
  XNOR2X4TS U1162 ( .A(n392), .B(n817), .Y(n827) );
  XNOR2X4TS U1163 ( .A(n393), .B(n818), .Y(n392) );
  AOI21X2TS U1164 ( .A0(n1812), .A1(n1810), .B0(n1449), .Y(n1820) );
  OAI2BB1X4TS U1165 ( .A0N(n1700), .A1N(sumOut[85]), .B0(n1699), .Y(n1701) );
  CLKINVX1TS U1166 ( .A(n1209), .Y(n1210) );
  NOR2X4TS U1167 ( .A(n842), .B(n1534), .Y(n1543) );
  NOR2X4TS U1168 ( .A(n1214), .B(n1205), .Y(n1221) );
  ADDFHX4TS U1169 ( .A(n1369), .B(n1368), .CI(n1367), .CO(n445), .S(n1370) );
  XOR2X2TS U1170 ( .A(n1377), .B(n1376), .Y(n395) );
  XOR2X1TS U1171 ( .A(n1821), .B(n1820), .Y(genblk1_0__mac_s[3]) );
  OAI2BB1X2TS U1172 ( .A0N(n723), .A1N(sumOut[65]), .B0(n725), .Y(n739) );
  OR2X2TS U1173 ( .A(n1237), .B(n1236), .Y(n396) );
  OAI21X2TS U1174 ( .A0(n652), .A1(n651), .B0(sumOut[27]), .Y(n650) );
  INVX2TS U1175 ( .A(n1009), .Y(n1013) );
  XOR2X4TS U1176 ( .A(n1047), .B(n1046), .Y(n1053) );
  NOR2BX2TS U1177 ( .AN(n130), .B(n1705), .Y(n831) );
  INVX2TS U1178 ( .A(n1829), .Y(n1830) );
  NAND2X2TS U1179 ( .A(n1613), .B(n1614), .Y(n1829) );
  NOR2X2TS U1180 ( .A(n644), .B(n645), .Y(n1296) );
  CLKINVX1TS U1181 ( .A(n1497), .Y(n400) );
  INVX2TS U1182 ( .A(n400), .Y(n401) );
  NAND2X4TS U1183 ( .A(n1583), .B(n1582), .Y(n1815) );
  NOR2X4TS U1184 ( .A(n1284), .B(n1078), .Y(n1090) );
  XOR2X4TS U1185 ( .A(n402), .B(n1015), .Y(n1038) );
  XOR2X4TS U1186 ( .A(n404), .B(n863), .Y(n866) );
  INVX2TS U1187 ( .A(n1275), .Y(n405) );
  NAND3X4TS U1188 ( .A(n453), .B(n452), .C(n454), .Y(n634) );
  OAI21X2TS U1189 ( .A0(n599), .A1(n598), .B0(n597), .Y(n653) );
  XOR2X4TS U1190 ( .A(n407), .B(n1679), .Y(n1698) );
  XOR2X4TS U1191 ( .A(n1683), .B(n1684), .Y(n407) );
  INVX2TS U1192 ( .A(n782), .Y(n785) );
  XNOR2X4TS U1193 ( .A(n826), .B(n792), .Y(n408) );
  NAND2X4TS U1194 ( .A(n1182), .B(n198), .Y(n1195) );
  XOR2X4TS U1195 ( .A(n626), .B(n627), .Y(n451) );
  OAI2BB1X2TS U1196 ( .A0N(n1595), .A1N(n1594), .B0(n1593), .Y(n1610) );
  XOR2X2TS U1197 ( .A(n455), .B(n461), .Y(n412) );
  OAI2BB1X4TS U1198 ( .A0N(n1217), .A1N(n1218), .B0(n1198), .Y(n414) );
  CLKAND2X2TS U1199 ( .A(n566), .B(n959), .Y(n1022) );
  XNOR2X4TS U1200 ( .A(n1245), .B(n1244), .Y(n1215) );
  OR2X4TS U1201 ( .A(n244), .B(n1499), .Y(n1246) );
  OAI2BB1X2TS U1202 ( .A0N(n1241), .A1N(sumOut[75]), .B0(n1240), .Y(n1256) );
  OR2X2TS U1203 ( .A(n1058), .B(n1057), .Y(n415) );
  NOR2X6TS U1204 ( .A(n1764), .B(n1763), .Y(n1770) );
  NAND2X4TS U1205 ( .A(n1782), .B(n1781), .Y(n1791) );
  OAI21X1TS U1206 ( .A0(n443), .A1(n1774), .B0(sumOut[87]), .Y(n1773) );
  OAI2BB1X4TS U1207 ( .A0N(n439), .A1N(n1120), .B0(n1119), .Y(n1121) );
  CLKINVX1TS U1208 ( .A(n1099), .Y(n1103) );
  NOR2X6TS U1209 ( .A(n1058), .B(n1057), .Y(n1280) );
  XOR2X2TS U1210 ( .A(n1125), .B(n1126), .Y(n1112) );
  XOR2X4TS U1211 ( .A(n1000), .B(n977), .Y(n984) );
  NAND2X4TS U1212 ( .A(n1329), .B(n1328), .Y(n1341) );
  NAND2X4TS U1213 ( .A(n1329), .B(n824), .Y(n1536) );
  NAND2X4TS U1214 ( .A(n1329), .B(n1111), .Y(n1127) );
  XOR2X4TS U1215 ( .A(n1179), .B(n1202), .Y(n418) );
  CLKINVX1TS U1216 ( .A(n1940), .Y(n419) );
  INVX2TS U1217 ( .A(n420), .Y(n421) );
  NAND2BX4TS U1218 ( .AN(n1364), .B(n1305), .Y(n1375) );
  INVX2TS U1219 ( .A(n1703), .Y(n422) );
  INVX2TS U1220 ( .A(n1788), .Y(n1703) );
  OAI21X2TS U1221 ( .A0(sumOut[85]), .A1(n1700), .B0(n1698), .Y(n1699) );
  XOR2X4TS U1222 ( .A(n885), .B(n884), .Y(n433) );
  NOR2BX4TS U1223 ( .AN(n199), .B(n1309), .Y(n1368) );
  CLKINVX1TS U1224 ( .A(n1883), .Y(n649) );
  NAND2X1TS U1225 ( .A(n1883), .B(n1887), .Y(n1889) );
  OAI2BB1X4TS U1226 ( .A0N(n689), .A1N(n688), .B0(n687), .Y(n728) );
  OAI2BB1X2TS U1227 ( .A0N(n1607), .A1N(n1608), .B0(n1606), .Y(n1614) );
  OAI21X1TS U1228 ( .A0(sumOut[65]), .A1(n723), .B0(n724), .Y(n725) );
  NOR2X8TS U1229 ( .A(n1262), .B(n506), .Y(n1106) );
  OAI21X2TS U1230 ( .A0(n996), .A1(n997), .B0(n994), .Y(n995) );
  OAI2BB1X4TS U1231 ( .A0N(n1663), .A1N(n1665), .B0(n1636), .Y(n1671) );
  OAI21X2TS U1232 ( .A0(n868), .A1(n869), .B0(n866), .Y(n867) );
  BUFX20TS U1233 ( .A(n1340), .Y(n1689) );
  INVX4TS U1234 ( .A(n1366), .Y(n425) );
  NOR2X4TS U1235 ( .A(n2059), .B(n2061), .Y(n1678) );
  XNOR2X4TS U1236 ( .A(n1655), .B(n1654), .Y(n1661) );
  NAND2X1TS U1237 ( .A(n1643), .B(n223), .Y(n1644) );
  ADDFHX2TS U1238 ( .A(n1428), .B(n1429), .CI(n1427), .S(n428) );
  ADDFHX2TS U1239 ( .A(n1428), .B(n1429), .CI(n1427), .CO(n1476), .S(n1451) );
  NOR2X4TS U1240 ( .A(n1362), .B(sumOut[33]), .Y(n1912) );
  OAI2BB1X4TS U1241 ( .A0N(n561), .A1N(n560), .B0(n595), .Y(n565) );
  NOR2X4TS U1242 ( .A(n1904), .B(n1804), .Y(n1403) );
  INVX2TS U1243 ( .A(n1904), .Y(n1905) );
  XOR2X4TS U1244 ( .A(n1697), .B(sumOut[85]), .Y(n1652) );
  INVX4TS U1245 ( .A(n193), .Y(n1647) );
  XOR2X1TS U1246 ( .A(n1083), .B(n1082), .Y(genblk1_4__mac_s[7]) );
  OAI2BB1X4TS U1247 ( .A0N(n1663), .A1N(n1665), .B0(n1636), .Y(n430) );
  NOR2X8TS U1248 ( .A(n1625), .B(n823), .Y(n1539) );
  OAI21X2TS U1249 ( .A0(n1398), .A1(n1397), .B0(sumOut[37]), .Y(n1396) );
  XOR2X4TS U1250 ( .A(n418), .B(n431), .Y(n434) );
  NAND2X4TS U1251 ( .A(n1388), .B(n1387), .Y(n1906) );
  NAND3BX2TS U1252 ( .AN(n1601), .B(n1827), .C(n1832), .Y(n1834) );
  NOR2X2TS U1253 ( .A(n1582), .B(n1583), .Y(n1601) );
  XNOR2X1TS U1254 ( .A(n1295), .B(n1294), .Y(genblk1_7__mac_s[5]) );
  OAI21X2TS U1255 ( .A0(n1222), .A1(n1221), .B0(n1224), .Y(n1197) );
  XOR2X2TS U1256 ( .A(n1041), .B(n1040), .Y(n1043) );
  XOR2X4TS U1257 ( .A(n434), .B(n414), .Y(n1235) );
  OAI2BB1X1TS U1258 ( .A0N(n1639), .A1N(n1629), .B0(n1638), .Y(n1627) );
  NAND2X2TS U1259 ( .A(n476), .B(n475), .Y(n477) );
  CLKINVX1TS U1260 ( .A(n1922), .Y(n435) );
  INVX2TS U1261 ( .A(n435), .Y(n436) );
  NAND2X4TS U1262 ( .A(n198), .B(n555), .Y(n573) );
  XOR2X4TS U1263 ( .A(n908), .B(n907), .Y(n437) );
  XOR2X4TS U1264 ( .A(n771), .B(n769), .Y(n773) );
  NAND2X1TS U1265 ( .A(n202), .B(n777), .Y(n770) );
  AND2X4TS U1266 ( .A(n807), .B(n806), .Y(n803) );
  OAI21X2TS U1267 ( .A0(n1266), .A1(n1267), .B0(n421), .Y(n1265) );
  ADDHX4TS U1268 ( .A(n610), .B(n274), .CO(n625), .S(n614) );
  NAND2X4TS U1269 ( .A(n565), .B(n564), .Y(n590) );
  NOR2X4TS U1270 ( .A(n1443), .B(n506), .Y(n475) );
  NAND2X4TS U1271 ( .A(n1061), .B(n1060), .Y(n1286) );
  OAI2BB1X4TS U1272 ( .A0N(sumOut[45]), .A1N(n1034), .B0(n972), .Y(n1060) );
  NOR2X4TS U1273 ( .A(n437), .B(n922), .Y(n1492) );
  CLKBUFX2TS U1274 ( .A(n237), .Y(n441) );
  INVX4TS U1275 ( .A(n889), .Y(n837) );
  AOI21X4TS U1276 ( .A0(n1866), .A1(n1864), .B0(n608), .Y(n1872) );
  XOR2X4TS U1277 ( .A(n1136), .B(n1137), .Y(n1113) );
  OAI2BB1X2TS U1278 ( .A0N(n443), .A1N(n1774), .B0(n1773), .Y(n1784) );
  XOR2X4TS U1279 ( .A(n1045), .B(n1044), .Y(n1047) );
  XOR2X4TS U1280 ( .A(n694), .B(n665), .Y(n666) );
  OAI2BB1X2TS U1281 ( .A0N(n1375), .A1N(sumOut[35]), .B0(n1317), .Y(n1387) );
  OAI21X2TS U1282 ( .A0(n2075), .A1(n181), .B0(n2072), .Y(n522) );
  OAI21X2TS U1283 ( .A0(n2080), .A1(n2083), .B0(n2081), .Y(n2069) );
  NOR2X2TS U1284 ( .A(sumOut[91]), .B(n468), .Y(n2080) );
  NOR2X4TS U1285 ( .A(n929), .B(n928), .Y(n442) );
  ADDFHX2TS U1286 ( .A(n1778), .B(n1777), .CI(n1776), .S(n443) );
  ADDFHX2TS U1287 ( .A(n1778), .B(n1777), .CI(n1776), .CO(n1797), .S(n1775) );
  OAI21X2TS U1288 ( .A0(n859), .A1(n858), .B0(n860), .Y(n845) );
  OAI21X1TS U1289 ( .A0(n1735), .A1(n1732), .B0(n1733), .Y(n1495) );
  NOR2X2TS U1290 ( .A(n1633), .B(n1348), .Y(n1354) );
  XOR2X1TS U1291 ( .A(n444), .B(n860), .Y(n447) );
  XOR2X4TS U1292 ( .A(n1380), .B(n445), .Y(n448) );
  NOR2X4TS U1293 ( .A(n1214), .B(n1301), .Y(n1359) );
  OAI21X4TS U1294 ( .A0(n1820), .A1(n1817), .B0(n1818), .Y(n1565) );
  NOR2X4TS U1295 ( .A(n1454), .B(sumOut[3]), .Y(n1817) );
  NAND2X2TS U1296 ( .A(n1454), .B(sumOut[3]), .Y(n1818) );
  NAND2X2TS U1297 ( .A(n623), .B(n621), .Y(n576) );
  XOR2X4TS U1298 ( .A(n1353), .B(n1373), .Y(n1362) );
  XOR2X4TS U1299 ( .A(n448), .B(n1378), .Y(n1382) );
  NAND2X4TS U1300 ( .A(n962), .B(n961), .Y(n1034) );
  NAND2X2TS U1301 ( .A(n1015), .B(n366), .Y(n962) );
  NAND2X2TS U1302 ( .A(n1365), .B(n1363), .Y(n1305) );
  XOR2X4TS U1303 ( .A(n1034), .B(n449), .Y(n1035) );
  OAI2BB1X2TS U1304 ( .A0N(n1498), .A1N(n401), .B0(n1496), .Y(n1507) );
  OAI21X2TS U1305 ( .A0(n1498), .A1(n401), .B0(sumOut[77]), .Y(n1496) );
  OAI2BB1X4TS U1306 ( .A0N(n1045), .A1N(n1044), .B0(n1031), .Y(n1042) );
  XOR2X4TS U1307 ( .A(n451), .B(n625), .Y(n619) );
  NAND2X4TS U1308 ( .A(n626), .B(n625), .Y(n452) );
  NAND2X2TS U1309 ( .A(n884), .B(n882), .Y(n857) );
  OAI21X4TS U1310 ( .A0(n1872), .A1(n1869), .B0(n1870), .Y(n643) );
  NAND2BX4TS U1311 ( .AN(n1204), .B(n1203), .Y(n1241) );
  NAND2X2TS U1312 ( .A(n1202), .B(n1201), .Y(n1203) );
  NAND2X2TS U1313 ( .A(n1460), .B(n1459), .Y(n1461) );
  NAND2X2TS U1314 ( .A(n1477), .B(n215), .Y(n1561) );
  OAI2BB1X4TS U1315 ( .A0N(sumOut[25]), .A1N(n635), .B0(n582), .Y(n644) );
  NOR2X4TS U1316 ( .A(n678), .B(n1181), .Y(n1226) );
  BUFX8TS U1317 ( .A(n1659), .Y(n678) );
  NOR2X4TS U1318 ( .A(n678), .B(n691), .Y(n705) );
  NAND2BX2TS U1319 ( .AN(n1645), .B(n1644), .Y(n1697) );
  OAI21X2TS U1320 ( .A0(n785), .A1(n786), .B0(n783), .Y(n784) );
  NAND2X2TS U1321 ( .A(n198), .B(n959), .Y(n1028) );
  OAI2BB1X2TS U1322 ( .A0N(n771), .A1N(n769), .B0(n768), .Y(n798) );
  NOR2X2TS U1323 ( .A(n765), .B(n1432), .Y(n806) );
  INVX2TS U1324 ( .A(sumOut[55]), .Y(n792) );
  OAI21X1TS U1325 ( .A0(n1170), .A1(n1171), .B0(sumOut[98]), .Y(n1169) );
  INVX2TS U1326 ( .A(n1003), .Y(n1006) );
  INVX2TS U1327 ( .A(sumOut[97]), .Y(n1133) );
  OAI21X1TS U1328 ( .A0(n1569), .A1(sumOut[5]), .B0(n1567), .Y(n1568) );
  XOR2X1TS U1329 ( .A(n1049), .B(n1048), .Y(n1052) );
  OAI2BB1X2TS U1330 ( .A0N(n1798), .A1N(n1797), .B0(n1796), .Y(n1799) );
  OAI21X1TS U1331 ( .A0(n1797), .A1(n1798), .B0(sumOut[88]), .Y(n1796) );
  NAND2X2TS U1332 ( .A(n1230), .B(sumOut[73]), .Y(n2029) );
  INVX2TS U1333 ( .A(n1990), .Y(n713) );
  AOI21X2TS U1334 ( .A0(n1931), .A1(n1933), .B0(n1054), .Y(n1946) );
  INVX2TS U1335 ( .A(n1126), .Y(n1129) );
  INVX2TS U1336 ( .A(n1150), .Y(n1111) );
  NAND2X2TS U1337 ( .A(n193), .B(n761), .Y(n819) );
  INVX2TS U1338 ( .A(n967), .Y(n980) );
  NAND2X2TS U1339 ( .A(n563), .B(n562), .Y(n564) );
  INVX2TS U1340 ( .A(n1007), .Y(n981) );
  INVX2TS U1341 ( .A(n1714), .Y(n824) );
  INVX2TS U1342 ( .A(n326), .Y(n668) );
  NAND2X1TS U1343 ( .A(n1123), .B(n968), .Y(n1009) );
  INVX2TS U1344 ( .A(n1014), .Y(n961) );
  NAND2X1TS U1345 ( .A(n566), .B(n260), .Y(n480) );
  AND2X4TS U1346 ( .A(n1657), .B(n1656), .Y(n1654) );
  INVX2TS U1347 ( .A(n1725), .Y(n1726) );
  INVX2TS U1348 ( .A(n1977), .Y(n1978) );
  AOI21X2TS U1349 ( .A0(n1091), .A1(n1095), .B0(n1066), .Y(n1067) );
  AOI21X2TS U1350 ( .A0(n1521), .A1(n1525), .B0(n1166), .Y(n1167) );
  INVX2TS U1351 ( .A(n1404), .Y(n1405) );
  CLKAND2X2TS U1352 ( .A(n2101), .B(genblk1_2__mac_biasesStored[9]), .Y(n464)
         );
  INVX2TS U1353 ( .A(n2044), .Y(n2060) );
  CLKBUFX2TS U1354 ( .A(n2094), .Y(n2113) );
  CLKBUFX2TS U1355 ( .A(n2112), .Y(n2101) );
  CLKBUFX2TS U1356 ( .A(n2110), .Y(n2123) );
  CLKBUFX2TS U1357 ( .A(n2127), .Y(n2118) );
  CLKBUFX2TS U1358 ( .A(n2094), .Y(n2115) );
  CLKBUFX2TS U1359 ( .A(n2111), .Y(n2114) );
  CLKBUFX2TS U1360 ( .A(n2112), .Y(n2117) );
  CLKBUFX2TS U1361 ( .A(n2110), .Y(n2122) );
  CLKBUFX2TS U1362 ( .A(n2111), .Y(n2124) );
  INVX2TS U1363 ( .A(n1832), .Y(n1615) );
  NAND2BXLTS U1364 ( .AN(genblk1_0__mac_biasesStored[9]), .B(n2118), .Y(n10)
         );
  NAND2BXLTS U1365 ( .AN(genblk1_7__mac_biasesStored[9]), .B(n2123), .Y(n94)
         );
  INVX2TS U1366 ( .A(n944), .Y(n757) );
  XNOR2X1TS U1367 ( .A(n1495), .B(n1494), .Y(genblk1_1__mac_s[5]) );
  NAND2BXLTS U1368 ( .AN(genblk1_2__mac_biasesStored[9]), .B(n2128), .Y(n540)
         );
  INVX2TS U1369 ( .A(n464), .Y(n2130) );
  NAND2BXLTS U1370 ( .AN(genblk1_8__mac_biasesStored[9]), .B(n2124), .Y(n106)
         );
  NAND2BXLTS U1371 ( .AN(genblk1_6__mac_biasesStored[9]), .B(n2128), .Y(n82)
         );
  NAND2BXLTS U1372 ( .AN(genblk1_4__mac_biasesStored[9]), .B(n2122), .Y(n543)
         );
  NAND2BXLTS U1373 ( .AN(genblk1_1__mac_biasesStored[9]), .B(n2114), .Y(n22)
         );
  AND2X4TS U1374 ( .A(n1486), .B(n1485), .Y(n1487) );
  NAND2BXLTS U1375 ( .AN(genblk1_3__mac_biasesStored[9]), .B(n2117), .Y(n548)
         );
  INVX2TS U1376 ( .A(n1520), .Y(n1523) );
  NAND2X1TS U1377 ( .A(n2095), .B(genblk1_9__mac_biasesStored[9]), .Y(n537) );
  NAND2X1TS U1378 ( .A(n2086), .B(n1528), .Y(n2088) );
  NAND2X1TS U1379 ( .A(n2099), .B(genblk1_7__mac_biasesStored[9]), .Y(n523) );
  NAND2BXLTS U1380 ( .AN(genblk1_5__mac_biasesStored[9]), .B(n2113), .Y(n70)
         );
  NAND2X1TS U1381 ( .A(n2104), .B(genblk1_5__mac_biasesStored[9]), .Y(n526) );
  NAND2X1TS U1382 ( .A(n2098), .B(genblk1_0__mac_biasesStored[9]), .Y(n531) );
  NAND2BXLTS U1383 ( .AN(genblk1_9__mac_biasesStored[9]), .B(n2115), .Y(n118)
         );
  OAI21X1TS U1384 ( .A0(n2027), .A1(n1290), .B0(n210), .Y(n1295) );
  NAND2X1TS U1385 ( .A(n2109), .B(genblk1_4__mac_biasesStored[9]), .Y(n528) );
  XNOR2X1TS U1386 ( .A(n1283), .B(n1282), .Y(genblk1_4__mac_s[5]) );
  NAND2BX2TS U1387 ( .AN(n1938), .B(n1936), .Y(n1279) );
  INVX2TS U1388 ( .A(n464), .Y(n2131) );
  XNOR2X1TS U1389 ( .A(n1480), .B(n1479), .Y(genblk1_0__mac_s[5]) );
  OAI21X2TS U1390 ( .A0(n1458), .A1(n1457), .B0(n1456), .Y(n1480) );
  XOR2X2TS U1391 ( .A(n1736), .B(n1735), .Y(genblk1_1__mac_s[4]) );
  INVX2TS U1392 ( .A(n1732), .Y(n1734) );
  XOR2XLTS U1393 ( .A(n2052), .B(n2051), .Y(genblk1_8__mac_s[3]) );
  XOR2XLTS U1394 ( .A(n2032), .B(n2031), .Y(genblk1_7__mac_s[3]) );
  XOR2XLTS U1395 ( .A(n2003), .B(n2002), .Y(genblk1_6__mac_s[3]) );
  XOR2XLTS U1396 ( .A(n1947), .B(n1946), .Y(genblk1_4__mac_s[3]) );
  XOR2XLTS U1397 ( .A(n1916), .B(n1915), .Y(genblk1_3__mac_s[3]) );
  XOR2XLTS U1398 ( .A(n1873), .B(n1872), .Y(genblk1_2__mac_s[3]) );
  XOR2XLTS U1399 ( .A(n1852), .B(n1851), .Y(genblk1_1__mac_s[3]) );
  XOR2XLTS U1400 ( .A(n1921), .B(n1920), .Y(genblk1_3__mac_s[1]) );
  XOR2XLTS U1401 ( .A(n1826), .B(n1825), .Y(genblk1_0__mac_s[1]) );
  INVX2TS U1402 ( .A(n1421), .Y(n1422) );
  INVX2TS U1403 ( .A(weightsIn[22]), .Y(n1312) );
  INVX2TS U1404 ( .A(weightsIn[43]), .Y(n1181) );
  INVX2TS U1405 ( .A(n260), .Y(n469) );
  INVX2TS U1406 ( .A(n1301), .Y(n1311) );
  INVX2TS U1407 ( .A(n765), .Y(n777) );
  INVX2TS U1408 ( .A(n838), .Y(n851) );
  INVX2TS U1409 ( .A(n1327), .Y(n1328) );
  INVX2TS U1410 ( .A(n602), .Y(n609) );
  INVX2TS U1411 ( .A(weightsIn[12]), .Y(n602) );
  AND2X4TS U1412 ( .A(n198), .B(n851), .Y(n862) );
  INVX2TS U1413 ( .A(n1346), .Y(n1351) );
  INVX2TS U1414 ( .A(n1626), .Y(n1621) );
  INVX6TS U1415 ( .A(n557), .Y(n595) );
  INVX4TS U1416 ( .A(n1316), .Y(n1376) );
  CLKINVX1TS U1417 ( .A(weightsIn[55]), .Y(n467) );
  NOR2X1TS U1418 ( .A(n469), .B(n188), .Y(n2070) );
  NAND2X1TS U1419 ( .A(sumOut[91]), .B(n468), .Y(n2081) );
  XOR2X4TS U1420 ( .A(n480), .B(n479), .Y(n476) );
  INVX2TS U1421 ( .A(weightsIn[56]), .Y(n506) );
  INVX2TS U1422 ( .A(n2066), .Y(n473) );
  CLKINVX1TS U1423 ( .A(weightsIn[57]), .Y(n505) );
  AND2X4TS U1424 ( .A(n489), .B(n1019), .Y(n487) );
  NOR2X4TS U1425 ( .A(n1417), .B(n506), .Y(n486) );
  XOR2X4TS U1426 ( .A(n487), .B(n486), .Y(n503) );
  NAND2X4TS U1427 ( .A(n482), .B(n483), .Y(n485) );
  NAND2X2TS U1428 ( .A(n484), .B(sumOut[93]), .Y(n2077) );
  NAND2X4TS U1429 ( .A(n487), .B(n486), .Y(n488) );
  NOR2X4TS U1430 ( .A(n1468), .B(n506), .Y(n510) );
  XOR2X4TS U1431 ( .A(n494), .B(n493), .Y(n511) );
  XOR2X4TS U1432 ( .A(n495), .B(n511), .Y(n516) );
  OAI2BB1X4TS U1433 ( .A0N(n503), .A1N(n502), .B0(n501), .Y(n514) );
  NAND2X4TS U1434 ( .A(n1152), .B(sumOut[94]), .Y(n1156) );
  INVX2TS U1435 ( .A(n1156), .Y(n504) );
  INVX2TS U1436 ( .A(n504), .Y(n2072) );
  NOR2X4TS U1437 ( .A(n1468), .B(n505), .Y(n1107) );
  XOR2X4TS U1438 ( .A(n1107), .B(n1106), .Y(n507) );
  XOR2X4TS U1439 ( .A(n507), .B(n1104), .Y(n1098) );
  INVX2TS U1440 ( .A(weightsIn[59]), .Y(n1150) );
  XOR2X4TS U1441 ( .A(n1118), .B(sumOut[95]), .Y(n513) );
  XOR2X4TS U1442 ( .A(n1115), .B(n513), .Y(n519) );
  NAND2X2TS U1443 ( .A(n518), .B(n519), .Y(n1154) );
  CLKINVX1TS U1444 ( .A(n1155), .Y(n520) );
  NAND2X1TS U1445 ( .A(n1154), .B(n520), .Y(n521) );
  CLKBUFX2TS U1446 ( .A(clr), .Y(n539) );
  CLKBUFX2TS U1447 ( .A(n539), .Y(n2091) );
  CLKBUFX2TS U1448 ( .A(n2091), .Y(n535) );
  CLKBUFX2TS U1449 ( .A(n535), .Y(n2099) );
  CLKBUFX2TS U1450 ( .A(n2091), .Y(n2108) );
  NAND2X1TS U1451 ( .A(n2108), .B(genblk1_6__mac_biasesStored[9]), .Y(n81) );
  CLKBUFX2TS U1452 ( .A(n2091), .Y(n2104) );
  CLKBUFX2TS U1453 ( .A(n535), .Y(n2109) );
  CLKBUFX2TS U1454 ( .A(n539), .Y(n2094) );
  CLKBUFX2TS U1455 ( .A(n2094), .Y(n2093) );
  CLKBUFX2TS U1456 ( .A(n2093), .Y(n2097) );
  CLKBUFX2TS U1457 ( .A(n2097), .Y(n2102) );
  NAND2X1TS U1458 ( .A(n2102), .B(genblk1_3__mac_biasesStored[9]), .Y(n45) );
  CLKBUFX2TS U1459 ( .A(n2097), .Y(n2098) );
  NAND2X1TS U1460 ( .A(n539), .B(genblk1_1__mac_biasesStored[9]), .Y(n533) );
  CLKBUFX2TS U1461 ( .A(n535), .Y(n2092) );
  CLKBUFX2TS U1462 ( .A(n2092), .Y(n2106) );
  NAND2X1TS U1463 ( .A(n2106), .B(genblk1_8__mac_biasesStored[9]), .Y(n105) );
  CLKBUFX2TS U1464 ( .A(n2092), .Y(n2095) );
  CLKBUFX2TS U1465 ( .A(n539), .Y(n2128) );
  CLKBUFX2TS U1466 ( .A(n2115), .Y(n2127) );
  CLKBUFX2TS U1467 ( .A(n2093), .Y(n2112) );
  CLKBUFX2TS U1468 ( .A(n2093), .Y(n2110) );
  CLKBUFX2TS U1469 ( .A(n2127), .Y(n2111) );
  CLKBUFX2TS U1470 ( .A(n82), .Y(n2132) );
  INVX2TS U1471 ( .A(weightsIn[17]), .Y(n656) );
  OR2X2TS U1472 ( .A(n1659), .B(n656), .Y(n577) );
  INVX2TS U1473 ( .A(n555), .Y(n567) );
  INVX2TS U1474 ( .A(weightsIn[16]), .Y(n593) );
  INVX2TS U1475 ( .A(weightsIn[14]), .Y(n604) );
  NAND2X4TS U1476 ( .A(n555), .B(n195), .Y(n561) );
  XNOR2X4TS U1477 ( .A(n560), .B(n561), .Y(n558) );
  INVX2TS U1478 ( .A(n593), .Y(n556) );
  AND2X4TS U1479 ( .A(n556), .B(n198), .Y(n557) );
  XNOR2X4TS U1480 ( .A(n558), .B(n595), .Y(n578) );
  OAI21X2TS U1481 ( .A0(n579), .A1(n577), .B0(n578), .Y(n559) );
  XOR2X4TS U1482 ( .A(n584), .B(sumOut[26]), .Y(n570) );
  INVX2TS U1483 ( .A(n560), .Y(n563) );
  INVX2TS U1484 ( .A(n561), .Y(n562) );
  NOR2X4TS U1485 ( .A(n1262), .B(n567), .Y(n596) );
  XOR2X4TS U1486 ( .A(n596), .B(n598), .Y(n568) );
  XOR2X4TS U1487 ( .A(n568), .B(n595), .Y(n586) );
  XOR2X4TS U1488 ( .A(n569), .B(n586), .Y(n585) );
  XOR2X4TS U1489 ( .A(n570), .B(n585), .Y(n645) );
  INVX2TS U1490 ( .A(n604), .Y(n572) );
  AND2X8TS U1491 ( .A(n267), .B(n611), .Y(n622) );
  XOR2X4TS U1492 ( .A(n575), .B(n574), .Y(n623) );
  NOR2X4TS U1493 ( .A(n1468), .B(n604), .Y(n621) );
  INVX2TS U1494 ( .A(n635), .Y(n581) );
  XOR2X4TS U1495 ( .A(n578), .B(n577), .Y(n580) );
  XOR2X4TS U1496 ( .A(n580), .B(n413), .Y(n637) );
  OAI2BB1X2TS U1497 ( .A0N(n584), .A1N(n585), .B0(n583), .Y(n646) );
  INVX2TS U1498 ( .A(n590), .Y(n587) );
  OAI2BB1X4TS U1499 ( .A0N(n588), .A1N(n587), .B0(n586), .Y(n589) );
  XNOR2X4TS U1500 ( .A(n600), .B(n652), .Y(n647) );
  NOR2X2TS U1501 ( .A(n1417), .B(n602), .Y(n605) );
  NOR2X1TS U1502 ( .A(sumOut[21]), .B(n603), .Y(n1874) );
  NOR2X1TS U1503 ( .A(n1633), .B(n602), .Y(n1867) );
  NAND2X1TS U1504 ( .A(sumOut[21]), .B(n603), .Y(n1875) );
  OR2X4TS U1505 ( .A(sumOut[22]), .B(n607), .Y(n1864) );
  NAND2X1TS U1506 ( .A(sumOut[22]), .B(n607), .Y(n1863) );
  INVX2TS U1507 ( .A(n1863), .Y(n608) );
  AND2X4TS U1508 ( .A(n204), .B(n609), .Y(n627) );
  CLKBUFX2TS U1509 ( .A(n267), .Y(n612) );
  XOR2X4TS U1510 ( .A(n612), .B(n125), .Y(n620) );
  XOR2X4TS U1511 ( .A(n619), .B(n620), .Y(n616) );
  XOR2X4TS U1512 ( .A(n616), .B(n618), .Y(n617) );
  NOR2X4TS U1513 ( .A(n617), .B(sumOut[23]), .Y(n1869) );
  NAND2X2TS U1514 ( .A(n617), .B(sumOut[23]), .Y(n1870) );
  XOR2X4TS U1515 ( .A(n622), .B(n621), .Y(n624) );
  XOR2X4TS U1516 ( .A(n624), .B(n623), .Y(n633) );
  XOR2X4TS U1517 ( .A(n633), .B(n634), .Y(n628) );
  XOR2X4TS U1518 ( .A(n629), .B(n628), .Y(n638) );
  NOR2X4TS U1519 ( .A(n638), .B(sumOut[24]), .Y(n1879) );
  OAI2BB1X4TS U1520 ( .A0N(n631), .A1N(n630), .B0(n629), .Y(n632) );
  OAI2BB1X4TS U1521 ( .A0N(n634), .A1N(n441), .B0(n632), .Y(n640) );
  XOR2X4TS U1522 ( .A(n637), .B(n636), .Y(n639) );
  NOR2X8TS U1523 ( .A(n640), .B(n639), .Y(n1085) );
  NOR2X4TS U1524 ( .A(n1879), .B(n1085), .Y(n642) );
  NAND2X4TS U1525 ( .A(n638), .B(sumOut[24]), .Y(n1084) );
  NAND2X2TS U1526 ( .A(n640), .B(n639), .Y(n1087) );
  OAI21X4TS U1527 ( .A0(n1084), .A1(n1085), .B0(n1087), .Y(n641) );
  AOI21X4TS U1528 ( .A0(n642), .A1(n643), .B0(n641), .Y(n1888) );
  NAND2X2TS U1529 ( .A(n647), .B(n646), .Y(n833) );
  OAI21X2TS U1530 ( .A0(n649), .A1(n1888), .B0(n648), .Y(n661) );
  OAI2BB1X2TS U1531 ( .A0N(n652), .A1N(n651), .B0(n650), .Y(n659) );
  OR2X4TS U1532 ( .A(n659), .B(n658), .Y(n1887) );
  XOR2X1TS U1533 ( .A(n661), .B(n660), .Y(genblk1_2__mac_s[8]) );
  INVX2TS U1534 ( .A(weightsIn[39]), .Y(n667) );
  INVX2TS U1535 ( .A(weightsIn[40]), .Y(n663) );
  NOR2X4TS U1536 ( .A(n1434), .B(n663), .Y(n686) );
  XOR2X4TS U1537 ( .A(n664), .B(n686), .Y(n694) );
  INVX2TS U1538 ( .A(weightsIn[38]), .Y(n691) );
  INVX2TS U1539 ( .A(weightsIn[36]), .Y(n703) );
  NOR2X4TS U1540 ( .A(n1418), .B(n703), .Y(n671) );
  XOR2X4TS U1541 ( .A(n671), .B(n670), .Y(n673) );
  XOR2X4TS U1542 ( .A(n673), .B(n672), .Y(n698) );
  XOR2X4TS U1543 ( .A(n677), .B(n676), .Y(n706) );
  NOR2X2TS U1544 ( .A(n1417), .B(n703), .Y(n702) );
  INVX2TS U1545 ( .A(n705), .Y(n679) );
  OAI2BB1X4TS U1546 ( .A0N(n705), .A1N(n706), .B0(n681), .Y(n699) );
  OAI21X4TS U1547 ( .A0(n208), .A1(n697), .B0(n699), .Y(n683) );
  NAND2X2TS U1548 ( .A(n208), .B(n697), .Y(n682) );
  XOR2X4TS U1549 ( .A(n717), .B(n716), .Y(n684) );
  OAI2BB1X4TS U1550 ( .A0N(n715), .A1N(n423), .B0(n685), .Y(n719) );
  INVX2TS U1551 ( .A(weightsIn[41]), .Y(n951) );
  XOR2X4TS U1552 ( .A(n728), .B(n690), .Y(n692) );
  NOR2X4TS U1553 ( .A(n1418), .B(n691), .Y(n733) );
  XNOR2X4TS U1554 ( .A(n692), .B(n726), .Y(n724) );
  NOR2X8TS U1555 ( .A(n720), .B(n719), .Y(n2011) );
  XOR2X4TS U1556 ( .A(n700), .B(n699), .Y(n714) );
  NOR2X2TS U1557 ( .A(n714), .B(sumOut[63]), .Y(n1999) );
  NOR2X1TS U1558 ( .A(sumOut[61]), .B(n704), .Y(n2004) );
  NAND2X1TS U1559 ( .A(sumOut[61]), .B(n704), .Y(n2005) );
  OAI21X2TS U1560 ( .A0(n2004), .A1(n2007), .B0(n2005), .Y(n1993) );
  XNOR2X4TS U1561 ( .A(n706), .B(n705), .Y(n709) );
  XOR2X4TS U1562 ( .A(n709), .B(n708), .Y(n712) );
  INVX2TS U1563 ( .A(n712), .Y(n711) );
  NAND2X2TS U1564 ( .A(sumOut[62]), .B(n712), .Y(n1990) );
  AOI21X2TS U1565 ( .A0(n1993), .A1(n1991), .B0(n713), .Y(n2002) );
  OAI21X2TS U1566 ( .A0(n1999), .A1(n2002), .B0(n2000), .Y(n1996) );
  XOR2X4TS U1567 ( .A(n717), .B(n716), .Y(n718) );
  NAND2X2TS U1568 ( .A(n720), .B(n719), .Y(n2013) );
  OAI21X4TS U1569 ( .A0(n398), .A1(n2011), .B0(n2013), .Y(n721) );
  AOI21X4TS U1570 ( .A0(n722), .A1(n1996), .B0(n721), .Y(n1744) );
  OAI21X2TS U1571 ( .A0(n728), .A1(n729), .B0(n726), .Y(n727) );
  OAI2BB1X4TS U1572 ( .A0N(n729), .A1N(n728), .B0(n727), .Y(n754) );
  XOR2X4TS U1573 ( .A(n754), .B(sumOut[66]), .Y(n738) );
  NOR2X2TS U1574 ( .A(n842), .B(n663), .Y(n743) );
  XOR2X4TS U1575 ( .A(n744), .B(n743), .Y(n737) );
  NOR2X4TS U1576 ( .A(n1016), .B(n734), .Y(n749) );
  XOR2X4TS U1577 ( .A(n749), .B(n750), .Y(n736) );
  NAND2X2TS U1578 ( .A(n1329), .B(n735), .Y(n746) );
  XOR2X4TS U1579 ( .A(n736), .B(n746), .Y(n741) );
  XOR2X4TS U1580 ( .A(n737), .B(n741), .Y(n753) );
  XOR2X4TS U1581 ( .A(n738), .B(n753), .Y(n740) );
  NOR2X2TS U1582 ( .A(n740), .B(n739), .Y(n1738) );
  OAI21X2TS U1583 ( .A0(n744), .A1(n743), .B0(n741), .Y(n742) );
  XOR2X4TS U1584 ( .A(n949), .B(sumOut[67]), .Y(n751) );
  NOR2X2TS U1585 ( .A(n1715), .B(n663), .Y(n954) );
  CLKINVX1TS U1586 ( .A(n749), .Y(n747) );
  OAI2BB1X2TS U1587 ( .A0N(n750), .A1N(n749), .B0(n748), .Y(n952) );
  XOR2X4TS U1588 ( .A(n751), .B(n950), .Y(n755) );
  OAI2BB1X4TS U1589 ( .A0N(n754), .A1N(n753), .B0(n752), .Y(n756) );
  CLKINVX3TS U1590 ( .A(n945), .Y(n1737) );
  NAND2X4TS U1591 ( .A(n756), .B(n755), .Y(n944) );
  NOR2X1TS U1592 ( .A(n757), .B(n945), .Y(n758) );
  XOR2X1TS U1593 ( .A(n759), .B(n758), .Y(genblk1_6__mac_s[7]) );
  AND2X4TS U1594 ( .A(n761), .B(n211), .Y(n774) );
  INVX2TS U1595 ( .A(n761), .Y(n775) );
  NOR2X8TS U1596 ( .A(n775), .B(n1689), .Y(n789) );
  XOR2X4TS U1597 ( .A(n791), .B(n789), .Y(n764) );
  INVX2TS U1598 ( .A(weightsIn[34]), .Y(n1534) );
  XOR2X4TS U1599 ( .A(n763), .B(n783), .Y(n790) );
  XOR2X4TS U1600 ( .A(n764), .B(n790), .Y(n797) );
  INVX2TS U1601 ( .A(weightsIn[30]), .Y(n765) );
  OAI21X1TS U1602 ( .A0(n769), .A1(n771), .B0(n772), .Y(n768) );
  XOR2X4TS U1603 ( .A(n797), .B(n798), .Y(n780) );
  XOR2X4TS U1604 ( .A(n773), .B(n772), .Y(n800) );
  XOR2X4TS U1605 ( .A(n455), .B(n461), .Y(n804) );
  INVX2TS U1606 ( .A(weightsIn[35]), .Y(n1714) );
  OR2X2TS U1607 ( .A(n898), .B(n1714), .Y(n818) );
  INVX2TS U1608 ( .A(n1534), .Y(n787) );
  OAI2BB1X4TS U1609 ( .A0N(n798), .A1N(n427), .B0(n796), .Y(n813) );
  NOR2X4TS U1610 ( .A(n1274), .B(n1971), .Y(n816) );
  NOR2X4TS U1611 ( .A(n811), .B(sumOut[53]), .Y(n1959) );
  XOR2X4TS U1612 ( .A(n805), .B(n412), .Y(n809) );
  OR2X4TS U1613 ( .A(sumOut[52]), .B(n809), .Y(n1954) );
  XOR2X1TS U1614 ( .A(n807), .B(n806), .Y(n808) );
  NOR2X1TS U1615 ( .A(sumOut[51]), .B(n808), .Y(n1964) );
  NOR2X1TS U1616 ( .A(n466), .B(n765), .Y(n1957) );
  NAND2X1TS U1617 ( .A(sumOut[50]), .B(n1957), .Y(n1967) );
  NAND2X1TS U1618 ( .A(sumOut[51]), .B(n808), .Y(n1965) );
  NAND2X1TS U1619 ( .A(sumOut[52]), .B(n809), .Y(n1953) );
  INVX2TS U1620 ( .A(n1953), .Y(n810) );
  AOI21X4TS U1621 ( .A0(n1954), .A1(n1956), .B0(n810), .Y(n1963) );
  NAND2X2TS U1622 ( .A(n811), .B(sumOut[53]), .Y(n1960) );
  OAI21X4TS U1623 ( .A0(n1959), .A1(n1963), .B0(n1960), .Y(n1277) );
  NAND2X4TS U1624 ( .A(n812), .B(sumOut[54]), .Y(n1969) );
  NAND2X2TS U1625 ( .A(n813), .B(n814), .Y(n1973) );
  OAI21X4TS U1626 ( .A0(n1969), .A1(n1971), .B0(n1973), .Y(n815) );
  XOR2X4TS U1627 ( .A(n1547), .B(sumOut[56]), .Y(n825) );
  INVX2TS U1628 ( .A(n819), .Y(n821) );
  XNOR2X1TS U1629 ( .A(n831), .B(n1982), .Y(genblk1_5__mac_s[6]) );
  CLKINVX1TS U1630 ( .A(n832), .Y(n834) );
  XOR2X1TS U1631 ( .A(n836), .B(n835), .Y(genblk1_2__mac_s[7]) );
  INVX2TS U1632 ( .A(weightsIn[7]), .Y(n889) );
  INVX2TS U1633 ( .A(weightsIn[10]), .Y(n838) );
  INVX2TS U1634 ( .A(weightsIn[9]), .Y(n886) );
  OAI21X2TS U1635 ( .A0(n854), .A1(n460), .B0(n855), .Y(n840) );
  INVX2TS U1636 ( .A(weightsIn[11]), .Y(n878) );
  NOR2X4TS U1637 ( .A(n745), .B(n886), .Y(n850) );
  XOR2X4TS U1638 ( .A(n850), .B(n848), .Y(n844) );
  OR2X4TS U1639 ( .A(n1619), .B(n838), .Y(n846) );
  XNOR2X4TS U1640 ( .A(n844), .B(n846), .Y(n860) );
  XOR2X4TS U1641 ( .A(n872), .B(sumOut[16]), .Y(n852) );
  OAI2BB1X4TS U1642 ( .A0N(n182), .A1N(n850), .B0(n849), .Y(n868) );
  NOR2X2TS U1643 ( .A(n134), .B(n838), .Y(n869) );
  XOR2X4TS U1644 ( .A(n852), .B(n873), .Y(n927) );
  XOR2X4TS U1645 ( .A(n460), .B(n854), .Y(n856) );
  XOR2X4TS U1646 ( .A(n856), .B(n855), .Y(n884) );
  NOR2X4TS U1647 ( .A(n926), .B(n927), .Y(n1858) );
  OR2X4TS U1648 ( .A(n1423), .B(n878), .Y(n880) );
  OAI2BB1X4TS U1649 ( .A0N(n865), .A1N(n862), .B0(n864), .Y(n879) );
  OAI2BB1X4TS U1650 ( .A0N(n869), .A1N(n868), .B0(n867), .Y(n875) );
  XOR2X4TS U1651 ( .A(n870), .B(n875), .Y(n929) );
  OAI21X4TS U1652 ( .A0(n209), .A1(n873), .B0(sumOut[16]), .Y(n871) );
  OAI2BB1X4TS U1653 ( .A0N(n209), .A1N(n873), .B0(n871), .Y(n928) );
  NOR2X4TS U1654 ( .A(n928), .B(n929), .Y(n1552) );
  NOR2X4TS U1655 ( .A(n1858), .B(n442), .Y(n1481) );
  OAI21X1TS U1656 ( .A0(n876), .A1(n875), .B0(sumOut[17]), .Y(n874) );
  OAI2BB1X1TS U1657 ( .A0N(n876), .A1N(n875), .B0(n874), .Y(n931) );
  OR2X2TS U1658 ( .A(n594), .B(n878), .Y(n936) );
  OR2X4TS U1659 ( .A(n931), .B(n930), .Y(n1486) );
  NAND2X2TS U1660 ( .A(n1481), .B(n1486), .Y(n934) );
  NOR2X4TS U1661 ( .A(n898), .B(n886), .Y(n894) );
  OAI2BB1X2TS U1662 ( .A0N(n890), .A1N(n888), .B0(n896), .Y(n891) );
  XOR2X4TS U1663 ( .A(n433), .B(n905), .Y(n903) );
  XOR2X4TS U1664 ( .A(n897), .B(n896), .Y(n910) );
  NOR2X2TS U1665 ( .A(n898), .B(n843), .Y(n916) );
  OAI2BB1X4TS U1666 ( .A0N(n905), .A1N(n433), .B0(n904), .Y(n922) );
  XOR2X4TS U1667 ( .A(n907), .B(n908), .Y(n923) );
  NOR2X1TS U1668 ( .A(n1051), .B(n887), .Y(n1846) );
  OAI21X2TS U1669 ( .A0(n1853), .A1(n1856), .B0(n1854), .Y(n1845) );
  NOR2X2TS U1670 ( .A(sumOut[12]), .B(n918), .Y(n917) );
  INVX2TS U1671 ( .A(n917), .Y(n1843) );
  INVX2TS U1672 ( .A(n1842), .Y(n919) );
  OAI21X4TS U1673 ( .A0(n1491), .A1(n1492), .B0(n1493), .Y(n924) );
  AOI21X4TS U1674 ( .A0(n925), .A1(n1489), .B0(n924), .Y(n1861) );
  NAND2X4TS U1675 ( .A(n927), .B(n926), .Y(n1860) );
  NAND2X2TS U1676 ( .A(n929), .B(n928), .Y(n1553) );
  OAI21X4TS U1677 ( .A0(n1860), .A1(n1552), .B0(n1553), .Y(n1482) );
  NAND2X1TS U1678 ( .A(n931), .B(n930), .Y(n1485) );
  INVX2TS U1679 ( .A(n1485), .Y(n932) );
  ADDFHX2TS U1680 ( .A(n936), .B(n935), .CI(sumOut[18]), .CO(n937), .S(n930)
         );
  INVX2TS U1681 ( .A(n937), .Y(n939) );
  NOR2X2TS U1682 ( .A(sumOut[19]), .B(n939), .Y(n938) );
  INVX2TS U1683 ( .A(n938), .Y(n941) );
  NAND2X1TS U1684 ( .A(sumOut[19]), .B(n939), .Y(n940) );
  AND2X2TS U1685 ( .A(n941), .B(n940), .Y(n942) );
  NAND2BX2TS U1686 ( .AN(n1738), .B(n1737), .Y(n947) );
  INVX2TS U1687 ( .A(n1742), .Y(n946) );
  OAI21X2TS U1688 ( .A0(n1744), .A1(n947), .B0(n946), .Y(n958) );
  OAI21X2TS U1689 ( .A0(n950), .A1(n949), .B0(sumOut[67]), .Y(n948) );
  OAI2BB1X2TS U1690 ( .A0N(n950), .A1N(n949), .B0(n948), .Y(n956) );
  ADDFHX2TS U1691 ( .A(n954), .B(n953), .CI(n952), .CO(n1745), .S(n950) );
  NAND2X1TS U1692 ( .A(n956), .B(n955), .Y(n1739) );
  NAND2XLTS U1693 ( .A(n1741), .B(n1739), .Y(n957) );
  XNOR2X1TS U1694 ( .A(n958), .B(n957), .Y(genblk1_6__mac_s[8]) );
  INVX2TS U1695 ( .A(n968), .Y(n990) );
  INVX2TS U1696 ( .A(weightsIn[25]), .Y(n1030) );
  XOR2X4TS U1697 ( .A(n964), .B(n963), .Y(n960) );
  INVX2TS U1698 ( .A(weightsIn[27]), .Y(n1017) );
  INVX2TS U1699 ( .A(weightsIn[26]), .Y(n1029) );
  OAI2BB1X2TS U1700 ( .A0N(n406), .A1N(n966), .B0(n965), .Y(n976) );
  INVX2TS U1701 ( .A(weightsIn[29]), .Y(n1007) );
  XOR2X4TS U1702 ( .A(n976), .B(n975), .Y(n971) );
  NAND2X1TS U1703 ( .A(n877), .B(n280), .Y(n967) );
  NAND2X4TS U1704 ( .A(n968), .B(n1691), .Y(n985) );
  XOR2X4TS U1705 ( .A(n971), .B(n973), .Y(n1036) );
  OAI2BB1X4TS U1706 ( .A0N(n975), .A1N(n976), .B0(n974), .Y(n1000) );
  OAI2BB1X4TS U1707 ( .A0N(n980), .A1N(n979), .B0(n978), .Y(n997) );
  INVX4TS U1708 ( .A(n1183), .Y(n1326) );
  XOR2X4TS U1709 ( .A(n997), .B(n996), .Y(n983) );
  XNOR2X4TS U1710 ( .A(n988), .B(n985), .Y(n982) );
  XOR2X4TS U1711 ( .A(n982), .B(n986), .Y(n994) );
  XOR2X4TS U1712 ( .A(n983), .B(n994), .Y(n1001) );
  XOR2X4TS U1713 ( .A(n984), .B(n1001), .Y(n1061) );
  INVX2TS U1714 ( .A(n985), .Y(n989) );
  OAI21X2TS U1715 ( .A0(n989), .A1(n988), .B0(n986), .Y(n987) );
  OR2X4TS U1716 ( .A(n1326), .B(n1007), .Y(n1012) );
  XOR2X4TS U1717 ( .A(n1013), .B(n1012), .Y(n992) );
  XOR2X4TS U1718 ( .A(n1002), .B(n993), .Y(n998) );
  OAI2BB1X2TS U1719 ( .A0N(n997), .A1N(n996), .B0(n995), .Y(n1003) );
  OAI21X2TS U1720 ( .A0(n1001), .A1(n1000), .B0(sumOut[46]), .Y(n999) );
  OR2X2TS U1721 ( .A(n594), .B(n1007), .Y(n1070) );
  INVX2TS U1722 ( .A(n1012), .Y(n1010) );
  OAI2BB1X2TS U1723 ( .A0N(n1010), .A1N(n1009), .B0(n1008), .Y(n1011) );
  OAI2BB1X2TS U1724 ( .A0N(n1013), .A1N(n1012), .B0(n1011), .Y(n1069) );
  OR2X4TS U1725 ( .A(n1065), .B(n1064), .Y(n1095) );
  NAND2X1TS U1726 ( .A(n1090), .B(n1095), .Y(n1068) );
  INVX2TS U1727 ( .A(weightsIn[24]), .Y(n1050) );
  INVX2TS U1728 ( .A(n1050), .Y(n1018) );
  NOR2X2TS U1729 ( .A(n1028), .B(n1027), .Y(n1024) );
  XOR2X4TS U1730 ( .A(n1038), .B(n1039), .Y(n1033) );
  XOR2X4TS U1731 ( .A(n1021), .B(n1022), .Y(n1040) );
  XOR2X4TS U1732 ( .A(n1028), .B(n235), .Y(n1045) );
  NOR2X2TS U1733 ( .A(n244), .B(n1030), .Y(n1048) );
  OAI21X2TS U1734 ( .A0(n1044), .A1(n1045), .B0(n1046), .Y(n1031) );
  OAI21X4TS U1735 ( .A0(n1040), .A1(n1041), .B0(n1042), .Y(n1032) );
  OAI2BB1X4TS U1736 ( .A0N(n1040), .A1N(n1041), .B0(n1032), .Y(n1037) );
  XOR2X4TS U1737 ( .A(n1033), .B(n1037), .Y(n1056) );
  NOR2X4TS U1738 ( .A(n1056), .B(sumOut[44]), .Y(n1938) );
  XOR2X4TS U1739 ( .A(n1036), .B(n1035), .Y(n1058) );
  NOR2X4TS U1740 ( .A(n1938), .B(n1280), .Y(n1059) );
  XOR2X4TS U1741 ( .A(n1043), .B(n1042), .Y(n1055) );
  NOR2X4TS U1742 ( .A(n1055), .B(sumOut[43]), .Y(n1943) );
  OR2X4TS U1743 ( .A(sumOut[42]), .B(n1053), .Y(n1931) );
  NOR2X1TS U1744 ( .A(n1051), .B(n1050), .Y(n1934) );
  NAND2X1TS U1745 ( .A(sumOut[41]), .B(n1052), .Y(n1949) );
  NAND2X1TS U1746 ( .A(n1053), .B(sumOut[42]), .Y(n1930) );
  NAND2X2TS U1747 ( .A(n1055), .B(sumOut[43]), .Y(n1945) );
  OAI21X4TS U1748 ( .A0(n1943), .A1(n1946), .B0(n1945), .Y(n1936) );
  NAND2X4TS U1749 ( .A(n1056), .B(sumOut[44]), .Y(n1937) );
  NAND2X2TS U1750 ( .A(n1058), .B(n1057), .Y(n1281) );
  NAND2X2TS U1751 ( .A(n1063), .B(n1062), .Y(n1079) );
  NAND2X1TS U1752 ( .A(n1065), .B(n1064), .Y(n1094) );
  OAI21X2TS U1753 ( .A0(n1068), .A1(n1287), .B0(n1067), .Y(n1077) );
  ADDFHX2TS U1754 ( .A(n1070), .B(n1069), .CI(sumOut[48]), .CO(n1071), .S(
        n1064) );
  INVX2TS U1755 ( .A(n1071), .Y(n1073) );
  NOR2X1TS U1756 ( .A(sumOut[49]), .B(n1073), .Y(n1072) );
  CLKINVX1TS U1757 ( .A(n1072), .Y(n1075) );
  NAND2X1TS U1758 ( .A(sumOut[49]), .B(n1073), .Y(n1074) );
  AND2X2TS U1759 ( .A(n1075), .B(n1074), .Y(n1076) );
  XOR2X1TS U1760 ( .A(n1077), .B(n1076), .Y(genblk1_4__mac_s[9]) );
  OAI21X2TS U1761 ( .A0(n410), .A1(n1287), .B0(n1286), .Y(n1083) );
  NAND2X1TS U1762 ( .A(n1080), .B(n1079), .Y(n1081) );
  OA21X4TS U1763 ( .A0(n1872), .A1(n1869), .B0(n1870), .Y(n1882) );
  CLKINVX1TS U1764 ( .A(n1085), .Y(n1086) );
  NAND2X1TS U1765 ( .A(n1087), .B(n1086), .Y(n1088) );
  INVX2TS U1766 ( .A(n1090), .Y(n1093) );
  INVX2TS U1767 ( .A(n1091), .Y(n1092) );
  OAI21X2TS U1768 ( .A0(n1093), .A1(n1287), .B0(n1092), .Y(n1097) );
  XOR2X1TS U1769 ( .A(n1097), .B(n1096), .Y(genblk1_4__mac_s[8]) );
  INVX2TS U1770 ( .A(n1102), .Y(n1100) );
  OAI2BB1X4TS U1771 ( .A0N(n1100), .A1N(n1099), .B0(n1098), .Y(n1101) );
  OAI2BB1X4TS U1772 ( .A0N(n1102), .A1N(n1103), .B0(n1101), .Y(n1122) );
  XOR2X4TS U1773 ( .A(n1122), .B(sumOut[96]), .Y(n1114) );
  OAI2BB1X2TS U1774 ( .A0N(n1107), .A1N(n1106), .B0(n1105), .Y(n1136) );
  INVX2TS U1775 ( .A(n1109), .Y(n1124) );
  NAND2X2TS U1776 ( .A(n491), .B(n1109), .Y(n1125) );
  NAND2X2TS U1777 ( .A(n194), .B(n1110), .Y(n1126) );
  XOR2X4TS U1778 ( .A(n1112), .B(n1127), .Y(n1134) );
  XOR2X4TS U1779 ( .A(n1113), .B(n1134), .Y(n1119) );
  XOR2X4TS U1780 ( .A(n1114), .B(n1119), .Y(n1161) );
  INVX2TS U1781 ( .A(n1118), .Y(n1116) );
  OAI2BB1X2TS U1782 ( .A0N(n1118), .A1N(sumOut[95]), .B0(n1117), .Y(n1160) );
  NOR2X2TS U1783 ( .A(n1161), .B(n1160), .Y(n2085) );
  CLKINVX1TS U1784 ( .A(n1122), .Y(n1120) );
  OAI2BB1X4TS U1785 ( .A0N(n1122), .A1N(sumOut[96]), .B0(n1121), .Y(n1163) );
  OR2X2TS U1786 ( .A(n1326), .B(n1150), .Y(n1149) );
  XOR2X4TS U1787 ( .A(n1149), .B(n1142), .Y(n1132) );
  NAND2X4TS U1788 ( .A(n1129), .B(n1128), .Y(n1143) );
  NAND2X4TS U1789 ( .A(n1145), .B(n1143), .Y(n1130) );
  NAND2BX4TS U1790 ( .AN(n1144), .B(n1130), .Y(n1131) );
  XOR2X4TS U1791 ( .A(n1132), .B(n1131), .Y(n1140) );
  XOR2X4TS U1792 ( .A(n1140), .B(n1133), .Y(n1138) );
  OAI21X2TS U1793 ( .A0(n1137), .A1(n1136), .B0(n1134), .Y(n1135) );
  XNOR2X4TS U1794 ( .A(n1138), .B(n1141), .Y(n1162) );
  INVX2TS U1795 ( .A(n1142), .Y(n1148) );
  OAI21X2TS U1796 ( .A0(n1145), .A1(n1144), .B0(n1143), .Y(n1146) );
  OAI21X2TS U1797 ( .A0(n1148), .A1(n1149), .B0(n1146), .Y(n1147) );
  OR2X2TS U1798 ( .A(n1625), .B(n1150), .Y(n1171) );
  NAND2X2TS U1799 ( .A(n1520), .B(n1525), .Y(n1168) );
  NOR2X4TS U1800 ( .A(n226), .B(sumOut[94]), .Y(n1153) );
  NOR2X4TS U1801 ( .A(n1153), .B(n1155), .Y(n1159) );
  AOI21X4TS U1802 ( .A0(n1158), .A1(n1159), .B0(n1157), .Y(n2087) );
  NAND2X1TS U1803 ( .A(n1165), .B(n1164), .Y(n1524) );
  OAI21X2TS U1804 ( .A0(n1168), .A1(n2087), .B0(n1167), .Y(n1176) );
  INVX2TS U1805 ( .A(n1172), .Y(n1173) );
  NAND2X1TS U1806 ( .A(sumOut[99]), .B(n1173), .Y(n1174) );
  INVX2TS U1807 ( .A(n254), .Y(n1205) );
  INVX2TS U1808 ( .A(weightsIn[46]), .Y(n1261) );
  INVX2TS U1809 ( .A(n1261), .Y(n1249) );
  BUFX4TS U1810 ( .A(weightsIn[45]), .Y(n1250) );
  XOR2X4TS U1811 ( .A(n1178), .B(n1212), .Y(n1202) );
  XOR2X4TS U1812 ( .A(n1179), .B(n1202), .Y(n1233) );
  INVX2TS U1813 ( .A(weightsIn[42]), .Y(n1180) );
  NOR2X4TS U1814 ( .A(n1647), .B(n1180), .Y(n1191) );
  INVX2TS U1815 ( .A(n1194), .Y(n1185) );
  OAI21X4TS U1816 ( .A0(n1190), .A1(n1191), .B0(n1192), .Y(n1187) );
  OAI2BB1X4TS U1817 ( .A0N(n1190), .A1N(n1191), .B0(n1187), .Y(n1231) );
  XOR2X4TS U1818 ( .A(n1189), .B(n1188), .Y(n1217) );
  XOR2X4TS U1819 ( .A(n1191), .B(n1190), .Y(n1193) );
  XOR2X4TS U1820 ( .A(n1193), .B(n1192), .Y(n1218) );
  XOR2X4TS U1821 ( .A(n1195), .B(n1194), .Y(n1222) );
  OAI2BB1X4TS U1822 ( .A0N(n1221), .A1N(n1222), .B0(n1197), .Y(n1219) );
  OAI21X4TS U1823 ( .A0(n1218), .A1(n1217), .B0(n1219), .Y(n1198) );
  OAI2BB1X4TS U1824 ( .A0N(n1231), .A1N(n418), .B0(n1200), .Y(n1237) );
  XOR2X4TS U1825 ( .A(n1241), .B(sumOut[75]), .Y(n1216) );
  CLKINVX1TS U1826 ( .A(weightsIn[45]), .Y(n1206) );
  NOR2X4TS U1827 ( .A(n1326), .B(n1206), .Y(n1254) );
  OR2X4TS U1828 ( .A(n1261), .B(n1302), .Y(n1253) );
  INVX2TS U1829 ( .A(weightsIn[47]), .Y(n1499) );
  XOR2X4TS U1830 ( .A(n1215), .B(n1242), .Y(n1239) );
  XOR2X4TS U1831 ( .A(n1216), .B(n1239), .Y(n1236) );
  XOR2X4TS U1832 ( .A(n1218), .B(n1217), .Y(n1220) );
  XOR2X4TS U1833 ( .A(n1220), .B(n1219), .Y(n1230) );
  XOR2X4TS U1834 ( .A(n1222), .B(n1221), .Y(n1223) );
  XOR2X4TS U1835 ( .A(n1224), .B(n1223), .Y(n1228) );
  OR2X4TS U1836 ( .A(sumOut[72]), .B(n1228), .Y(n2017) );
  NOR2X2TS U1837 ( .A(sumOut[71]), .B(n1227), .Y(n2033) );
  NAND2X1TS U1838 ( .A(sumOut[71]), .B(n1227), .Y(n2034) );
  OAI21X1TS U1839 ( .A0(n2033), .A1(n2036), .B0(n2034), .Y(n2019) );
  INVX2TS U1840 ( .A(n2016), .Y(n1229) );
  AOI21X4TS U1841 ( .A0(n2017), .A1(n2019), .B0(n1229), .Y(n2031) );
  OAI21X4TS U1842 ( .A0(n2028), .A1(n2031), .B0(n2029), .Y(n1289) );
  NAND2X4TS U1843 ( .A(n1235), .B(sumOut[74]), .Y(n1291) );
  NAND2X2TS U1844 ( .A(n1236), .B(n1237), .Y(n1293) );
  OAI21X1TS U1845 ( .A0(sumOut[75]), .A1(n1241), .B0(n1239), .Y(n1240) );
  NOR2X2TS U1846 ( .A(n842), .B(n1261), .Y(n1267) );
  XOR2X4TS U1847 ( .A(n1264), .B(n1267), .Y(n1255) );
  XOR2X4TS U1848 ( .A(n1255), .B(n1266), .Y(n1260) );
  OR2X4TS U1849 ( .A(n745), .B(n1499), .Y(n1502) );
  NOR2X4TS U1850 ( .A(n1261), .B(n1262), .Y(n1503) );
  XOR2X4TS U1851 ( .A(n1502), .B(n1503), .Y(n1263) );
  XOR2X4TS U1852 ( .A(n1500), .B(n1263), .Y(n1497) );
  XOR2X4TS U1853 ( .A(n1497), .B(sumOut[77]), .Y(n1268) );
  OAI2BB1X2TS U1854 ( .A0N(n1267), .A1N(n1266), .B0(n1265), .Y(n1498) );
  XOR2X4TS U1855 ( .A(n1498), .B(n1268), .Y(n1269) );
  NAND2X2TS U1856 ( .A(n1270), .B(n1269), .Y(n1504) );
  CLKINVX1TS U1857 ( .A(n1504), .Y(n1271) );
  NOR2X1TS U1858 ( .A(n1271), .B(n1505), .Y(n1272) );
  CLKINVX1TS U1859 ( .A(n1969), .Y(n1276) );
  INVX2TS U1860 ( .A(n1274), .Y(n1275) );
  NAND2BX2TS U1861 ( .AN(n1276), .B(n1275), .Y(n1278) );
  INVX2TS U1862 ( .A(n1277), .Y(n1970) );
  NAND2X1TS U1863 ( .A(n1281), .B(n415), .Y(n1282) );
  NAND2X1TS U1864 ( .A(n1286), .B(n1285), .Y(n1288) );
  XOR2X1TS U1865 ( .A(n1288), .B(n1287), .Y(genblk1_4__mac_s[6]) );
  INVX2TS U1866 ( .A(n1289), .Y(n2027) );
  INVX2TS U1867 ( .A(n1290), .Y(n2025) );
  NAND2X1TS U1868 ( .A(n1293), .B(n396), .Y(n1294) );
  CLKINVX1TS U1869 ( .A(n1296), .Y(n1297) );
  NAND2X1TS U1870 ( .A(n1298), .B(n1297), .Y(n1299) );
  XOR2X1TS U1871 ( .A(n1299), .B(n1888), .Y(genblk1_2__mac_s[6]) );
  INVX2TS U1872 ( .A(n250), .Y(n1348) );
  INVX2TS U1873 ( .A(weightsIn[20]), .Y(n1301) );
  INVX2TS U1874 ( .A(n262), .Y(n1309) );
  XOR2X4TS U1875 ( .A(n1304), .B(n1307), .Y(n1365) );
  NOR2X4TS U1876 ( .A(n1423), .B(n1301), .Y(n1363) );
  INVX2TS U1877 ( .A(weightsIn[23]), .Y(n1327) );
  XOR2X4TS U1878 ( .A(n1325), .B(n1322), .Y(n1314) );
  OAI2BB1X4TS U1879 ( .A0N(n1321), .A1N(n1320), .B0(n1319), .Y(n1336) );
  XOR2X4TS U1880 ( .A(n1336), .B(sumOut[36]), .Y(n1331) );
  XNOR2X4TS U1881 ( .A(n1331), .B(n1332), .Y(n1388) );
  OAI2BB1X4TS U1882 ( .A0N(n1333), .A1N(n1332), .B0(sumOut[36]), .Y(n1334) );
  XOR2X4TS U1883 ( .A(n1397), .B(sumOut[37]), .Y(n1345) );
  OR2X4TS U1884 ( .A(n842), .B(n1327), .Y(n1394) );
  XOR2X4TS U1885 ( .A(n1345), .B(n1398), .Y(n1390) );
  INVX2TS U1886 ( .A(weightsIn[18]), .Y(n1346) );
  XOR2X4TS U1887 ( .A(n1370), .B(n1372), .Y(n1353) );
  NOR2X4TS U1888 ( .A(n1417), .B(n1346), .Y(n1355) );
  NOR2X1TS U1889 ( .A(n1051), .B(n1346), .Y(n1902) );
  NAND2X1TS U1890 ( .A(sumOut[31]), .B(n1356), .Y(n1918) );
  INVX2TS U1891 ( .A(n1898), .Y(n1361) );
  NAND2X2TS U1892 ( .A(n1362), .B(sumOut[33]), .Y(n1914) );
  NOR2X4TS U1893 ( .A(n1382), .B(sumOut[34]), .Y(n1923) );
  XOR2X4TS U1894 ( .A(n1375), .B(n1374), .Y(n1377) );
  XOR2X4TS U1895 ( .A(n1377), .B(n1376), .Y(n1383) );
  OAI2BB1X4TS U1896 ( .A0N(n445), .A1N(n1380), .B0(n1379), .Y(n1384) );
  NAND2X4TS U1897 ( .A(n1382), .B(sumOut[34]), .Y(n1922) );
  NAND2X2TS U1898 ( .A(n1389), .B(n1390), .Y(n1806) );
  INVX2TS U1899 ( .A(n1407), .Y(n1391) );
  OAI21X2TS U1900 ( .A0(n1392), .A1(n1907), .B0(n1391), .Y(n1402) );
  OR2X2TS U1901 ( .A(n1647), .B(n1327), .Y(n1411) );
  OR2X4TS U1902 ( .A(n1399), .B(n1400), .Y(n1406) );
  NAND2X1TS U1903 ( .A(n1400), .B(n1399), .Y(n1404) );
  XOR2X1TS U1904 ( .A(n1402), .B(n1401), .Y(genblk1_3__mac_s[8]) );
  OAI21X2TS U1905 ( .A0(n1409), .A1(n1907), .B0(n1408), .Y(n1416) );
  INVX2TS U1906 ( .A(n1412), .Y(n1413) );
  NAND2X1TS U1907 ( .A(sumOut[39]), .B(n1413), .Y(n1414) );
  AND2X2TS U1908 ( .A(n272), .B(n1414), .Y(n1415) );
  XOR2X1TS U1909 ( .A(n1416), .B(n1415), .Y(genblk1_3__mac_s[9]) );
  INVX2TS U1910 ( .A(weightsIn[3]), .Y(n1577) );
  INVX2TS U1911 ( .A(n1426), .Y(n1433) );
  INVX2TS U1912 ( .A(weightsIn[4]), .Y(n1591) );
  XOR2X4TS U1913 ( .A(n1419), .B(n1463), .Y(n1460) );
  INVX2TS U1914 ( .A(weightsIn[2]), .Y(n1421) );
  NOR2X4TS U1915 ( .A(n1423), .B(n1421), .Y(n1459) );
  XOR2X4TS U1916 ( .A(n1460), .B(n1424), .Y(n1475) );
  XOR2X4TS U1917 ( .A(n1475), .B(n1476), .Y(n1436) );
  NOR2X2TS U1918 ( .A(n1434), .B(n1433), .Y(n1440) );
  XOR2X4TS U1919 ( .A(n1436), .B(n1473), .Y(n1437) );
  INVX2TS U1920 ( .A(n1457), .Y(n1439) );
  NAND2X4TS U1921 ( .A(n1437), .B(sumOut[4]), .Y(n1562) );
  CLKINVX1TS U1922 ( .A(n1562), .Y(n1438) );
  INVX2TS U1923 ( .A(n1438), .Y(n1456) );
  NAND2X2TS U1924 ( .A(n1439), .B(n1456), .Y(n1455) );
  NOR2X1TS U1925 ( .A(sumOut[1]), .B(n1444), .Y(n1822) );
  NOR2X1TS U1926 ( .A(n1051), .B(n1442), .Y(n1813) );
  NAND2X1TS U1927 ( .A(sumOut[0]), .B(n1813), .Y(n1825) );
  NAND2X1TS U1928 ( .A(sumOut[1]), .B(n1444), .Y(n1823) );
  OAI21X1TS U1929 ( .A0(n1822), .A1(n1825), .B0(n1823), .Y(n1812) );
  OR2X4TS U1930 ( .A(sumOut[2]), .B(n1448), .Y(n1810) );
  XOR2X4TS U1931 ( .A(n1453), .B(n1452), .Y(n1454) );
  INVX2TS U1932 ( .A(n1565), .Y(n1458) );
  XOR2X2TS U1933 ( .A(n1455), .B(n1458), .Y(genblk1_0__mac_s[4]) );
  OAI2BB1X4TS U1934 ( .A0N(n1466), .A1N(n1465), .B0(n1464), .Y(n1572) );
  INVX2TS U1935 ( .A(weightsIn[5]), .Y(n1609) );
  OR2X2TS U1936 ( .A(n1651), .B(n1609), .Y(n1573) );
  XOR2X4TS U1937 ( .A(n1572), .B(n1467), .Y(n1471) );
  INVX2TS U1938 ( .A(n1591), .Y(n1470) );
  XNOR2X4TS U1939 ( .A(n1471), .B(n1570), .Y(n1567) );
  XOR2X4TS U1940 ( .A(n1472), .B(n1567), .Y(n1477) );
  OAI2BB1X4TS U1941 ( .A0N(n1476), .A1N(n217), .B0(n1474), .Y(n1478) );
  NAND2X1TS U1942 ( .A(n1561), .B(n216), .Y(n1479) );
  INVX2TS U1943 ( .A(n1481), .Y(n1484) );
  INVX2TS U1944 ( .A(n1482), .Y(n1483) );
  OAI21X2TS U1945 ( .A0(n1861), .A1(n1484), .B0(n1483), .Y(n1488) );
  INVX2TS U1946 ( .A(n1489), .Y(n1735) );
  NAND2X1TS U1947 ( .A(n1493), .B(n450), .Y(n1494) );
  OAI2BB1X2TS U1948 ( .A0N(n1503), .A1N(n1502), .B0(n1501), .Y(n1511) );
  OR2X4TS U1949 ( .A(n1507), .B(n1506), .Y(n1729) );
  NAND2X2TS U1950 ( .A(n1724), .B(n1729), .Y(n1510) );
  OAI21X4TS U1951 ( .A0(n2022), .A1(n1505), .B0(n1504), .Y(n1725) );
  NAND2X1TS U1952 ( .A(n1507), .B(n1506), .Y(n1728) );
  ADDFHX2TS U1953 ( .A(n1512), .B(n1511), .CI(sumOut[78]), .CO(n1513), .S(
        n1506) );
  INVX2TS U1954 ( .A(n1513), .Y(n1515) );
  INVX2TS U1955 ( .A(n1514), .Y(n1517) );
  NAND2X1TS U1956 ( .A(sumOut[79]), .B(n1515), .Y(n1516) );
  NAND2X1TS U1957 ( .A(n1517), .B(n1516), .Y(n1518) );
  INVX2TS U1958 ( .A(n1521), .Y(n1522) );
  AND2X2TS U1959 ( .A(n1531), .B(n1530), .Y(n1532) );
  NOR2X2TS U1960 ( .A(n1647), .B(n1534), .Y(n1719) );
  OR2X8TS U1961 ( .A(n383), .B(n1714), .Y(n1718) );
  XNOR2X4TS U1962 ( .A(n1719), .B(n1718), .Y(n1540) );
  INVX2TS U1963 ( .A(n1535), .Y(n1538) );
  OAI2BB1X4TS U1964 ( .A0N(n1539), .A1N(n1538), .B0(n1537), .Y(n1716) );
  XNOR2X4TS U1965 ( .A(n1540), .B(n1716), .Y(n1713) );
  XOR2X4TS U1966 ( .A(n1713), .B(sumOut[57]), .Y(n1544) );
  XOR2X4TS U1967 ( .A(n1544), .B(n1712), .Y(n1548) );
  OAI2BB1X4TS U1968 ( .A0N(n394), .A1N(n1547), .B0(n1545), .Y(n1549) );
  NAND2X2TS U1969 ( .A(n1548), .B(n1549), .Y(n1706) );
  OAI21X2TS U1970 ( .A0(n1861), .A1(n1858), .B0(n1860), .Y(n1556) );
  INVX2TS U1971 ( .A(n442), .Y(n1554) );
  CLKINVX1TS U1972 ( .A(n1738), .Y(n1557) );
  NAND2X1TS U1973 ( .A(n1558), .B(n1557), .Y(n1559) );
  XOR2X1TS U1974 ( .A(n1559), .B(n1744), .Y(genblk1_6__mac_s[6]) );
  NOR2X4TS U1975 ( .A(n1560), .B(n1563), .Y(n1566) );
  OAI2BB1X2TS U1976 ( .A0N(sumOut[5]), .A1N(n1569), .B0(n1568), .Y(n1582) );
  OAI2BB1X4TS U1977 ( .A0N(n1573), .A1N(n1572), .B0(n1571), .Y(n1585) );
  XOR2X4TS U1978 ( .A(n1585), .B(sumOut[6]), .Y(n1581) );
  XOR2X4TS U1979 ( .A(n1594), .B(n1578), .Y(n1579) );
  OR2X4TS U1980 ( .A(n1619), .B(n1609), .Y(n1592) );
  XNOR2X4TS U1981 ( .A(n1579), .B(n1592), .Y(n1587) );
  XNOR2X4TS U1982 ( .A(n1580), .B(n1587), .Y(n1586) );
  XOR2X4TS U1983 ( .A(n1581), .B(n1586), .Y(n1583) );
  OAI2BB1X4TS U1984 ( .A0N(n1590), .A1N(n1589), .B0(n1588), .Y(n1608) );
  XOR2X4TS U1985 ( .A(n1608), .B(sumOut[7]), .Y(n1596) );
  OR2X2TS U1986 ( .A(n842), .B(n1609), .Y(n1611) );
  XOR2X4TS U1987 ( .A(n1596), .B(n1607), .Y(n1598) );
  NAND2X2TS U1988 ( .A(n1597), .B(n1598), .Y(n1602) );
  XOR2X1TS U1989 ( .A(n1600), .B(n1599), .Y(genblk1_0__mac_s[7]) );
  INVX2TS U1990 ( .A(n1601), .Y(n1828) );
  OR2X2TS U1991 ( .A(n1418), .B(n1609), .Y(n1836) );
  NOR2BX1TS U1992 ( .AN(n1829), .B(n1615), .Y(n1616) );
  INVX2TS U1993 ( .A(weightsIn[49]), .Y(n1626) );
  INVX2TS U1994 ( .A(weightsIn[50]), .Y(n1646) );
  INVX2TS U1995 ( .A(weightsIn[51]), .Y(n1692) );
  XNOR2X4TS U1996 ( .A(n1624), .B(n1643), .Y(n1640) );
  INVX2TS U1997 ( .A(weightsIn[48]), .Y(n1658) );
  XOR2X4TS U1998 ( .A(n1640), .B(n1627), .Y(n1669) );
  XOR2X4TS U1999 ( .A(n1630), .B(n458), .Y(n1665) );
  NOR2X2TS U2000 ( .A(n1635), .B(n1658), .Y(n1657) );
  OAI21X4TS U2001 ( .A0(n1665), .A1(n1663), .B0(n1666), .Y(n1636) );
  XOR2X4TS U2002 ( .A(n1669), .B(n430), .Y(n1637) );
  OAI21X4TS U2003 ( .A0(n1674), .A1(n1673), .B0(n1671), .Y(n1641) );
  OAI21X4TS U2004 ( .A0(n397), .A1(n1650), .B0(n1648), .Y(n1649) );
  OAI2BB1X4TS U2005 ( .A0N(n397), .A1N(n1650), .B0(n1649), .Y(n1683) );
  INVX2TS U2006 ( .A(weightsIn[53]), .Y(n1779) );
  OR2X2TS U2007 ( .A(n1651), .B(n1779), .Y(n1684) );
  XOR2X4TS U2008 ( .A(n1653), .B(n1634), .Y(n1655) );
  OR2X4TS U2009 ( .A(sumOut[82]), .B(n1661), .Y(n2039) );
  XOR2X1TS U2010 ( .A(n1657), .B(n1656), .Y(n1660) );
  NOR2X1TS U2011 ( .A(sumOut[81]), .B(n1660), .Y(n2053) );
  NAND2X1TS U2012 ( .A(sumOut[81]), .B(n1660), .Y(n2054) );
  OAI21X1TS U2013 ( .A0(n2053), .A1(n2056), .B0(n2054), .Y(n2041) );
  INVX2TS U2014 ( .A(n2038), .Y(n1662) );
  XOR2X4TS U2015 ( .A(n1665), .B(n1664), .Y(n1667) );
  XNOR2X4TS U2016 ( .A(n1667), .B(n1666), .Y(n1668) );
  NOR2X4TS U2017 ( .A(n1668), .B(sumOut[83]), .Y(n2048) );
  NAND2X2TS U2018 ( .A(n1668), .B(sumOut[83]), .Y(n2049) );
  OAI21X4TS U2019 ( .A0(n2051), .A1(n2048), .B0(n2049), .Y(n2044) );
  XOR2X4TS U2020 ( .A(n1669), .B(n430), .Y(n1670) );
  NAND2X4TS U2021 ( .A(n1670), .B(sumOut[84]), .Y(n2045) );
  OAI2BB1X2TS U2022 ( .A0N(n1673), .A1N(n1674), .B0(n1672), .Y(n1675) );
  NAND2X2TS U2023 ( .A(n1676), .B(n1675), .Y(n2063) );
  AOI21X4TS U2024 ( .A0(n1678), .A1(n2044), .B0(n1677), .Y(n1794) );
  OAI2BB1X4TS U2025 ( .A0N(n1684), .A1N(n1683), .B0(n1682), .Y(n1754) );
  XOR2X4TS U2026 ( .A(n1754), .B(sumOut[86]), .Y(n1696) );
  OAI2BB1X4TS U2027 ( .A0N(n1688), .A1N(n1687), .B0(n1686), .Y(n1757) );
  XOR2X4TS U2028 ( .A(n1696), .B(n1753), .Y(n1702) );
  NOR2X2TS U2029 ( .A(n1702), .B(n1701), .Y(n1788) );
  NAND2X1TS U2030 ( .A(n1703), .B(n1769), .Y(n1704) );
  XOR2X1TS U2031 ( .A(n1704), .B(n1794), .Y(genblk1_8__mac_s[6]) );
  NOR2X4TS U2032 ( .A(n1705), .B(n1708), .Y(n1976) );
  INVX2TS U2033 ( .A(n1976), .Y(n1710) );
  OAI21X4TS U2034 ( .A0(n1708), .A1(n1707), .B0(n1706), .Y(n1980) );
  INVX2TS U2035 ( .A(n1980), .Y(n1709) );
  OAI2BB1X4TS U2036 ( .A0N(n1719), .A1N(n1718), .B0(n1717), .Y(n1984) );
  OR2X4TS U2037 ( .A(n1721), .B(n1720), .Y(n1979) );
  XOR2X1TS U2038 ( .A(n1723), .B(n1722), .Y(genblk1_5__mac_s[8]) );
  NAND2X2TS U2039 ( .A(n1734), .B(n1733), .Y(n1736) );
  NAND3BX2TS U2040 ( .AN(n1738), .B(n1737), .C(n1741), .Y(n1743) );
  INVX2TS U2041 ( .A(n1739), .Y(n1740) );
  ADDFHX2TS U2042 ( .A(n1746), .B(sumOut[68]), .CI(n1745), .CO(n1747), .S(n955) );
  INVX2TS U2043 ( .A(n1747), .Y(n1748) );
  NAND2X1TS U2044 ( .A(sumOut[69]), .B(n1748), .Y(n1749) );
  OAI21X2TS U2045 ( .A0(n1794), .A1(n422), .B0(n1769), .Y(n1767) );
  OAI2BB1X4TS U2046 ( .A0N(n1754), .A1N(n1753), .B0(n1752), .Y(n1763) );
  OAI2BB1X4TS U2047 ( .A0N(n1758), .A1N(n1757), .B0(n1756), .Y(n1774) );
  XOR2X4TS U2048 ( .A(n1774), .B(sumOut[87]), .Y(n1762) );
  NOR2X2TS U2049 ( .A(n1418), .B(n243), .Y(n1778) );
  OR2X4TS U2050 ( .A(n134), .B(n1779), .Y(n1777) );
  XOR2X4TS U2051 ( .A(n1762), .B(n1775), .Y(n1764) );
  NAND2X2TS U2052 ( .A(n1764), .B(n1763), .Y(n1768) );
  NAND2X1TS U2053 ( .A(n1768), .B(n1787), .Y(n1765) );
  NAND2BX2TS U2054 ( .AN(n1788), .B(n1787), .Y(n1772) );
  INVX2TS U2055 ( .A(n1792), .Y(n1771) );
  NAND2X2TS U2056 ( .A(n1784), .B(n1783), .Y(n1789) );
  NAND3BX2TS U2057 ( .AN(n1788), .B(n1787), .C(n1791), .Y(n1795) );
  INVX2TS U2058 ( .A(n1789), .Y(n1790) );
  INVX2TS U2059 ( .A(n1799), .Y(n1800) );
  NAND2X1TS U2060 ( .A(sumOut[89]), .B(n1800), .Y(n1801) );
  NAND2X1TS U2061 ( .A(n268), .B(n1801), .Y(n1802) );
  OAI21X2TS U2062 ( .A0(n1907), .A1(n1904), .B0(n1906), .Y(n1808) );
  INVX2TS U2063 ( .A(n1804), .Y(n1805) );
  NAND2X1TS U2064 ( .A(n1810), .B(n1809), .Y(n1811) );
  XNOR2X1TS U2065 ( .A(n1812), .B(n1811), .Y(genblk1_0__mac_s[2]) );
  OR2X2TS U2066 ( .A(sumOut[0]), .B(n1813), .Y(n1814) );
  XOR2X1TS U2067 ( .A(n1816), .B(n1833), .Y(genblk1_0__mac_s[6]) );
  NAND2X1TS U2068 ( .A(n1819), .B(n1818), .Y(n1821) );
  INVX2TS U2069 ( .A(n1837), .Y(n1838) );
  NAND2X1TS U2070 ( .A(sumOut[9]), .B(n1838), .Y(n1839) );
  AND2X2TS U2071 ( .A(n273), .B(n1839), .Y(n1840) );
  NAND2X1TS U2072 ( .A(n1843), .B(n1842), .Y(n1844) );
  XNOR2X1TS U2073 ( .A(n1845), .B(n1844), .Y(genblk1_1__mac_s[2]) );
  OR2X2TS U2074 ( .A(sumOut[10]), .B(n1846), .Y(n1847) );
  CLKINVX1TS U2075 ( .A(n1848), .Y(n1849) );
  NAND2X1TS U2076 ( .A(n1850), .B(n1849), .Y(n1852) );
  CLKINVX1TS U2077 ( .A(n1858), .Y(n1859) );
  NAND2X1TS U2078 ( .A(n1860), .B(n1859), .Y(n1862) );
  XOR2X1TS U2079 ( .A(n1862), .B(n1861), .Y(genblk1_1__mac_s[6]) );
  NAND2X1TS U2080 ( .A(n1864), .B(n1863), .Y(n1865) );
  XNOR2X1TS U2081 ( .A(n1866), .B(n1865), .Y(genblk1_2__mac_s[2]) );
  OR2X2TS U2082 ( .A(sumOut[20]), .B(n1867), .Y(n1868) );
  CLKINVX1TS U2083 ( .A(n1869), .Y(n1871) );
  NAND2X1TS U2084 ( .A(n1871), .B(n1870), .Y(n1873) );
  INVX2TS U2085 ( .A(n1879), .Y(n1880) );
  XOR2X1TS U2086 ( .A(n1882), .B(n1881), .Y(genblk1_2__mac_s[4]) );
  INVX2TS U2087 ( .A(n1893), .Y(n1894) );
  NAND2X1TS U2088 ( .A(sumOut[29]), .B(n1894), .Y(n1895) );
  AND2X2TS U2089 ( .A(n270), .B(n1895), .Y(n1896) );
  NAND2X1TS U2090 ( .A(n1899), .B(n1898), .Y(n1900) );
  XNOR2X1TS U2091 ( .A(n1901), .B(n1900), .Y(genblk1_3__mac_s[2]) );
  OR2X2TS U2092 ( .A(sumOut[30]), .B(n1902), .Y(n1903) );
  NAND2X1TS U2093 ( .A(n1906), .B(n1905), .Y(n1908) );
  XOR2X1TS U2094 ( .A(n1908), .B(n1907), .Y(genblk1_3__mac_s[6]) );
  INVX2TS U2095 ( .A(n1909), .Y(n1924) );
  CLKINVX1TS U2096 ( .A(n1923), .Y(n1910) );
  NAND2X1TS U2097 ( .A(n436), .B(n1910), .Y(n1911) );
  XOR2X1TS U2098 ( .A(n1924), .B(n1911), .Y(genblk1_3__mac_s[4]) );
  CLKINVX1TS U2099 ( .A(n1912), .Y(n1913) );
  NAND2X1TS U2100 ( .A(n1914), .B(n1913), .Y(n1916) );
  OAI21X1TS U2101 ( .A0(n1924), .A1(n1923), .B0(n436), .Y(n1929) );
  NAND2X1TS U2102 ( .A(n1927), .B(n1926), .Y(n1928) );
  XNOR2X1TS U2103 ( .A(n1929), .B(n1928), .Y(genblk1_3__mac_s[5]) );
  NAND2X1TS U2104 ( .A(n1931), .B(n1930), .Y(n1932) );
  XNOR2X1TS U2105 ( .A(n1933), .B(n1932), .Y(genblk1_4__mac_s[2]) );
  OR2X2TS U2106 ( .A(sumOut[40]), .B(n1934), .Y(n1935) );
  CLKINVX1TS U2107 ( .A(n1937), .Y(n1940) );
  CLKINVX1TS U2108 ( .A(n1938), .Y(n1939) );
  NAND2BX2TS U2109 ( .AN(n1940), .B(n1939), .Y(n1941) );
  XOR2X1TS U2110 ( .A(n1942), .B(n1941), .Y(genblk1_4__mac_s[4]) );
  NAND2X1TS U2111 ( .A(n1945), .B(n1944), .Y(n1947) );
  NAND2X1TS U2112 ( .A(n1954), .B(n1953), .Y(n1955) );
  XNOR2X1TS U2113 ( .A(n1956), .B(n1955), .Y(genblk1_5__mac_s[2]) );
  OR2X2TS U2114 ( .A(sumOut[50]), .B(n1957), .Y(n1958) );
  NAND2X1TS U2115 ( .A(n1961), .B(n1960), .Y(n1962) );
  XOR2X1TS U2116 ( .A(n1962), .B(n1963), .Y(genblk1_5__mac_s[3]) );
  CLKINVX1TS U2117 ( .A(n1964), .Y(n1966) );
  CLKINVX1TS U2118 ( .A(n1971), .Y(n1972) );
  NAND2X1TS U2119 ( .A(n1973), .B(n1972), .Y(n1974) );
  XNOR2X1TS U2120 ( .A(n1975), .B(n1974), .Y(genblk1_5__mac_s[5]) );
  NAND2X2TS U2121 ( .A(n1976), .B(n1979), .Y(n1983) );
  AOI21X4TS U2122 ( .A0(n1980), .A1(n1979), .B0(n1978), .Y(n1981) );
  ADDFHX2TS U2123 ( .A(n1985), .B(n1984), .CI(sumOut[58]), .CO(n1986), .S(
        n1720) );
  INVX2TS U2124 ( .A(n1986), .Y(n1987) );
  NAND2X1TS U2125 ( .A(sumOut[59]), .B(n1987), .Y(n1988) );
  AND2X2TS U2126 ( .A(n275), .B(n1988), .Y(n1989) );
  NAND2X1TS U2127 ( .A(n1991), .B(n1990), .Y(n1992) );
  XNOR2X1TS U2128 ( .A(n1992), .B(n1993), .Y(genblk1_6__mac_s[2]) );
  OR2X2TS U2129 ( .A(sumOut[60]), .B(n1994), .Y(n1995) );
  INVX2TS U2130 ( .A(n1996), .Y(n2010) );
  XOR2X1TS U2131 ( .A(n2010), .B(n1998), .Y(genblk1_6__mac_s[4]) );
  CLKINVX1TS U2132 ( .A(n1999), .Y(n2001) );
  NAND2X1TS U2133 ( .A(n2000), .B(n2001), .Y(n2003) );
  OAI21X1TS U2134 ( .A0(n2010), .A1(n2009), .B0(n206), .Y(n2015) );
  CLKINVX1TS U2135 ( .A(n2011), .Y(n2012) );
  NAND2X1TS U2136 ( .A(n2013), .B(n2012), .Y(n2014) );
  XNOR2X1TS U2137 ( .A(n2015), .B(n2014), .Y(genblk1_6__mac_s[5]) );
  NAND2X1TS U2138 ( .A(n2017), .B(n2016), .Y(n2018) );
  XNOR2X1TS U2139 ( .A(n2019), .B(n2018), .Y(genblk1_7__mac_s[2]) );
  NAND2X1TS U2140 ( .A(n2025), .B(n210), .Y(n2026) );
  XOR2X1TS U2141 ( .A(n2027), .B(n2026), .Y(genblk1_7__mac_s[4]) );
  CLKINVX1TS U2142 ( .A(n2028), .Y(n2030) );
  NAND2X1TS U2143 ( .A(n2030), .B(n2029), .Y(n2032) );
  NAND2XLTS U2144 ( .A(n2035), .B(n2034), .Y(n2037) );
  NAND2X1TS U2145 ( .A(n2039), .B(n2038), .Y(n2040) );
  XNOR2X1TS U2146 ( .A(n2041), .B(n2040), .Y(genblk1_8__mac_s[2]) );
  OR2X2TS U2147 ( .A(sumOut[80]), .B(n2042), .Y(n2043) );
  AND2X2TS U2148 ( .A(n2043), .B(n2056), .Y(genblk1_8__mac_s[0]) );
  CLKBUFX2TS U2149 ( .A(n2045), .Y(n2058) );
  CLKINVX1TS U2150 ( .A(n2059), .Y(n2046) );
  XOR2X1TS U2151 ( .A(n2060), .B(n2047), .Y(genblk1_8__mac_s[4]) );
  INVX2TS U2152 ( .A(n2048), .Y(n2050) );
  NAND2X1TS U2153 ( .A(n2050), .B(n2049), .Y(n2052) );
  OAI21X1TS U2154 ( .A0(n2060), .A1(n2059), .B0(n2058), .Y(n2065) );
  NAND2X1TS U2155 ( .A(n2063), .B(n2062), .Y(n2064) );
  XNOR2X1TS U2156 ( .A(n2065), .B(n2064), .Y(genblk1_8__mac_s[5]) );
  NAND2X1TS U2157 ( .A(n2066), .B(n2067), .Y(n2068) );
  XNOR2X1TS U2158 ( .A(n2069), .B(n2068), .Y(genblk1_9__mac_s[2]) );
  OR2X2TS U2159 ( .A(sumOut[90]), .B(n2070), .Y(n2071) );
  XOR2X1TS U2160 ( .A(n2075), .B(n2074), .Y(genblk1_9__mac_s[4]) );
  NAND2X1TS U2161 ( .A(n180), .B(n2077), .Y(n2079) );
  XOR2X1TS U2162 ( .A(n2079), .B(n2078), .Y(genblk1_9__mac_s[3]) );
  XOR2X1TS U2163 ( .A(n2088), .B(n2087), .Y(genblk1_9__mac_s[6]) );
  CLKBUFX2TS U2164 ( .A(biasWriteEnable), .Y(n2129) );
  CLKBUFX2TS U2165 ( .A(n2129), .Y(n2089) );
  CLKBUFX2TS U2166 ( .A(n2089), .Y(n2135) );
  CLKBUFX2TS U2167 ( .A(n2089), .Y(n2134) );
  CLKBUFX2TS U2168 ( .A(n2089), .Y(n2137) );
  CLKBUFX2TS U2169 ( .A(n2089), .Y(n2090) );
  CLKBUFX2TS U2170 ( .A(n2090), .Y(n2139) );
  CLKBUFX2TS U2171 ( .A(n2090), .Y(n2140) );
  CLKBUFX2TS U2172 ( .A(n2090), .Y(n2141) );
  CLKBUFX2TS U2173 ( .A(n2090), .Y(n2142) );
  CLKBUFX2TS U2174 ( .A(n2129), .Y(n2133) );
  CLKBUFX2TS U2175 ( .A(biasWriteEnable), .Y(n2146) );
  CLKBUFX2TS U2176 ( .A(biasWriteEnable), .Y(n2147) );
  CLKBUFX2TS U2177 ( .A(n2097), .Y(n2107) );
  NAND2X1TS U2178 ( .A(n2107), .B(genblk1_3__mac_biasesStored[1]), .Y(n37) );
  NAND2X1TS U2179 ( .A(n2104), .B(genblk1_4__mac_biasesStored[1]), .Y(n49) );
  NAND2X1TS U2180 ( .A(n2102), .B(genblk1_2__mac_biasesStored[1]), .Y(n25) );
  NAND2X1TS U2181 ( .A(n2110), .B(genblk1_1__mac_biasesStored[1]), .Y(n13) );
  CLKBUFX2TS U2182 ( .A(n2092), .Y(n2103) );
  NAND2X1TS U2183 ( .A(n2103), .B(genblk1_5__mac_biasesStored[1]), .Y(n61) );
  NAND2X1TS U2184 ( .A(n2098), .B(genblk1_0__mac_biasesStored[1]), .Y(n1) );
  CLKBUFX2TS U2185 ( .A(n2091), .Y(n2096) );
  NAND2X1TS U2186 ( .A(n2096), .B(genblk1_7__mac_biasesStored[0]), .Y(n95) );
  NAND2X1TS U2187 ( .A(n2099), .B(genblk1_6__mac_biasesStored[1]), .Y(n73) );
  NAND2X1TS U2188 ( .A(n2099), .B(genblk1_6__mac_biasesStored[0]), .Y(n83) );
  NAND2X1TS U2189 ( .A(n2096), .B(genblk1_7__mac_biasesStored[1]), .Y(n85) );
  NAND2X1TS U2190 ( .A(n2107), .B(genblk1_3__mac_biasesStored[0]), .Y(n47) );
  NAND2X1TS U2191 ( .A(n2102), .B(genblk1_2__mac_biasesStored[0]), .Y(n35) );
  NAND2X1TS U2192 ( .A(n2095), .B(genblk1_8__mac_biasesStored[1]), .Y(n97) );
  NAND2X1TS U2193 ( .A(n2101), .B(genblk1_1__mac_biasesStored[0]), .Y(n23) );
  CLKBUFX2TS U2194 ( .A(n2092), .Y(n2105) );
  NAND2X1TS U2195 ( .A(n2105), .B(genblk1_9__mac_biasesStored[1]), .Y(n109) );
  CLKBUFX2TS U2196 ( .A(n2093), .Y(n2100) );
  NAND2X1TS U2197 ( .A(n2100), .B(genblk1_0__mac_biasesStored[0]), .Y(n11) );
  NAND2X1TS U2198 ( .A(n2100), .B(genblk1_0__mac_biasesStored[2]), .Y(n3) );
  NAND2X1TS U2199 ( .A(n2108), .B(genblk1_6__mac_biasesStored[2]), .Y(n75) );
  NAND2X1TS U2200 ( .A(n2094), .B(genblk1_1__mac_biasesStored[4]), .Y(n19) );
  NAND2X1TS U2201 ( .A(n2101), .B(genblk1_2__mac_biasesStored[4]), .Y(n31) );
  NAND2X1TS U2202 ( .A(n2095), .B(genblk1_8__mac_biasesStored[0]), .Y(n107) );
  NAND2X1TS U2203 ( .A(n2108), .B(genblk1_6__mac_biasesStored[4]), .Y(n79) );
  NAND2X1TS U2204 ( .A(n2103), .B(genblk1_5__mac_biasesStored[3]), .Y(n65) );
  NAND2X1TS U2205 ( .A(n2100), .B(genblk1_0__mac_biasesStored[3]), .Y(n5) );
  NAND2X1TS U2206 ( .A(n2096), .B(genblk1_7__mac_biasesStored[3]), .Y(n89) );
  NAND2X1TS U2207 ( .A(n2095), .B(genblk1_9__mac_biasesStored[4]), .Y(n115) );
  NAND2X1TS U2208 ( .A(n2105), .B(genblk1_9__mac_biasesStored[3]), .Y(n113) );
  NAND2X1TS U2209 ( .A(n2109), .B(genblk1_4__mac_biasesStored[4]), .Y(n55) );
  NAND2X1TS U2210 ( .A(n2096), .B(genblk1_7__mac_biasesStored[2]), .Y(n87) );
  NAND2X1TS U2211 ( .A(n2106), .B(genblk1_8__mac_biasesStored[4]), .Y(n103) );
  NAND2X1TS U2212 ( .A(n2098), .B(genblk1_1__mac_biasesStored[2]), .Y(n15) );
  NAND2X1TS U2213 ( .A(n2097), .B(genblk1_1__mac_biasesStored[3]), .Y(n17) );
  NAND2X1TS U2214 ( .A(n2098), .B(genblk1_3__mac_biasesStored[4]), .Y(n43) );
  NAND2X1TS U2215 ( .A(n2099), .B(genblk1_7__mac_biasesStored[4]), .Y(n91) );
  NAND2X1TS U2216 ( .A(n2104), .B(genblk1_4__mac_biasesStored[0]), .Y(n59) );
  NAND2X1TS U2217 ( .A(n2107), .B(genblk1_3__mac_biasesStored[3]), .Y(n41) );
  NAND2X1TS U2218 ( .A(n2100), .B(genblk1_0__mac_biasesStored[4]), .Y(n7) );
  NAND2X1TS U2219 ( .A(n2101), .B(genblk1_2__mac_biasesStored[3]), .Y(n29) );
  NAND2X1TS U2220 ( .A(n2103), .B(genblk1_5__mac_biasesStored[0]), .Y(n71) );
  NAND2X1TS U2221 ( .A(n2102), .B(genblk1_2__mac_biasesStored[2]), .Y(n27) );
  NAND2X1TS U2222 ( .A(n2103), .B(genblk1_5__mac_biasesStored[2]), .Y(n63) );
  NAND2X1TS U2223 ( .A(n2104), .B(genblk1_5__mac_biasesStored[4]), .Y(n67) );
  NAND2X1TS U2224 ( .A(n2105), .B(genblk1_9__mac_biasesStored[0]), .Y(n119) );
  NAND2X1TS U2225 ( .A(n2106), .B(genblk1_8__mac_biasesStored[2]), .Y(n99) );
  NAND2X1TS U2226 ( .A(n2105), .B(genblk1_9__mac_biasesStored[2]), .Y(n111) );
  NAND2X1TS U2227 ( .A(n2106), .B(genblk1_8__mac_biasesStored[3]), .Y(n101) );
  NAND2X1TS U2228 ( .A(n2107), .B(genblk1_3__mac_biasesStored[2]), .Y(n39) );
  NAND2X1TS U2229 ( .A(n2109), .B(genblk1_4__mac_biasesStored[3]), .Y(n53) );
  NAND2X1TS U2230 ( .A(n2108), .B(genblk1_6__mac_biasesStored[3]), .Y(n77) );
  NAND2X1TS U2231 ( .A(n2109), .B(genblk1_4__mac_biasesStored[2]), .Y(n51) );
  NAND2BXLTS U2232 ( .AN(genblk1_3__mac_biasesStored[4]), .B(n2117), .Y(n44)
         );
  NAND2BXLTS U2233 ( .AN(genblk1_7__mac_biasesStored[4]), .B(n2123), .Y(n92)
         );
  CLKBUFX2TS U2234 ( .A(n2127), .Y(n2116) );
  NAND2BXLTS U2235 ( .AN(genblk1_9__mac_biasesStored[4]), .B(n2116), .Y(n116)
         );
  NAND2BXLTS U2236 ( .AN(genblk1_8__mac_biasesStored[4]), .B(n2124), .Y(n104)
         );
  NAND2BXLTS U2237 ( .AN(genblk1_5__mac_biasesStored[4]), .B(n2113), .Y(n68)
         );
  NAND2BXLTS U2238 ( .AN(genblk1_7__mac_biasesStored[1]), .B(n2114), .Y(n86)
         );
  NAND2BXLTS U2239 ( .AN(genblk1_1__mac_biasesStored[2]), .B(n2122), .Y(n16)
         );
  NAND2BXLTS U2240 ( .AN(genblk1_2__mac_biasesStored[3]), .B(n2113), .Y(n30)
         );
  NAND2BXLTS U2241 ( .AN(genblk1_9__mac_biasesStored[3]), .B(n2116), .Y(n114)
         );
  NAND2BXLTS U2242 ( .AN(genblk1_0__mac_biasesStored[3]), .B(n2116), .Y(n6) );
  NAND2BXLTS U2243 ( .AN(genblk1_3__mac_biasesStored[2]), .B(n2117), .Y(n40)
         );
  CLKBUFX2TS U2244 ( .A(n2110), .Y(n2120) );
  NAND2BXLTS U2245 ( .AN(genblk1_6__mac_biasesStored[4]), .B(n2120), .Y(n80)
         );
  CLKBUFX2TS U2246 ( .A(n2111), .Y(n2119) );
  NAND2BXLTS U2247 ( .AN(genblk1_2__mac_biasesStored[4]), .B(n2119), .Y(n32)
         );
  CLKBUFX2TS U2248 ( .A(n2111), .Y(n2121) );
  NAND2BXLTS U2249 ( .AN(genblk1_8__mac_biasesStored[3]), .B(n2121), .Y(n102)
         );
  NAND2BXLTS U2250 ( .AN(genblk1_9__mac_biasesStored[1]), .B(n2118), .Y(n110)
         );
  NAND2BXLTS U2251 ( .AN(genblk1_5__mac_biasesStored[1]), .B(n2119), .Y(n62)
         );
  CLKBUFX2TS U2252 ( .A(n2112), .Y(n2125) );
  NAND2BXLTS U2253 ( .AN(genblk1_3__mac_biasesStored[3]), .B(n2125), .Y(n42)
         );
  NAND2BXLTS U2254 ( .AN(genblk1_8__mac_biasesStored[2]), .B(n2121), .Y(n100)
         );
  NAND2BXLTS U2255 ( .AN(genblk1_4__mac_biasesStored[4]), .B(n2125), .Y(n56)
         );
  NAND2BXLTS U2256 ( .AN(genblk1_7__mac_biasesStored[3]), .B(n2121), .Y(n90)
         );
  NAND2BXLTS U2257 ( .AN(genblk1_1__mac_biasesStored[3]), .B(n2123), .Y(n18)
         );
  NAND2BXLTS U2258 ( .AN(genblk1_4__mac_biasesStored[2]), .B(clr), .Y(n52) );
  NAND2BXLTS U2259 ( .AN(genblk1_7__mac_biasesStored[2]), .B(n2114), .Y(n88)
         );
  NAND2BXLTS U2260 ( .AN(genblk1_9__mac_biasesStored[2]), .B(n2118), .Y(n112)
         );
  NAND2BXLTS U2261 ( .AN(genblk1_8__mac_biasesStored[1]), .B(n2115), .Y(n98)
         );
  NAND2BXLTS U2262 ( .AN(genblk1_6__mac_biasesStored[3]), .B(n2120), .Y(n78)
         );
  NAND2BXLTS U2263 ( .AN(genblk1_4__mac_biasesStored[1]), .B(clr), .Y(n50) );
  NAND2BXLTS U2264 ( .AN(genblk1_2__mac_biasesStored[2]), .B(n535), .Y(n28) );
  NAND2BXLTS U2265 ( .AN(genblk1_4__mac_biasesStored[3]), .B(n2113), .Y(n54)
         );
  NAND2BXLTS U2266 ( .AN(genblk1_6__mac_biasesStored[2]), .B(n2120), .Y(n76)
         );
  NAND2BXLTS U2267 ( .AN(genblk1_1__mac_biasesStored[4]), .B(n2114), .Y(n20)
         );
  NAND2BXLTS U2268 ( .AN(genblk1_0__mac_biasesStored[2]), .B(n2115), .Y(n4) );
  NAND2BXLTS U2269 ( .AN(genblk1_0__mac_biasesStored[4]), .B(n2116), .Y(n8) );
  NAND2BXLTS U2270 ( .AN(genblk1_5__mac_biasesStored[3]), .B(n2119), .Y(n66)
         );
  NAND2BXLTS U2271 ( .AN(genblk1_6__mac_biasesStored[1]), .B(n2122), .Y(n74)
         );
  NAND2BXLTS U2272 ( .AN(genblk1_3__mac_biasesStored[1]), .B(n2117), .Y(n38)
         );
  NAND2BXLTS U2273 ( .AN(genblk1_9__mac_biasesStored[0]), .B(n2118), .Y(n120)
         );
  NAND2BXLTS U2274 ( .AN(genblk1_5__mac_biasesStored[2]), .B(n2119), .Y(n64)
         );
  NAND2BXLTS U2275 ( .AN(genblk1_2__mac_biasesStored[1]), .B(n2112), .Y(n26)
         );
  NAND2BXLTS U2276 ( .AN(genblk1_1__mac_biasesStored[1]), .B(n2120), .Y(n14)
         );
  NAND2BXLTS U2277 ( .AN(genblk1_0__mac_biasesStored[1]), .B(n2121), .Y(n2) );
  NAND2BXLTS U2278 ( .AN(genblk1_7__mac_biasesStored[0]), .B(n2124), .Y(n96)
         );
  NAND2BXLTS U2279 ( .AN(genblk1_6__mac_biasesStored[0]), .B(n2122), .Y(n84)
         );
  NAND2BXLTS U2280 ( .AN(genblk1_1__mac_biasesStored[0]), .B(n2123), .Y(n24)
         );
  NAND2BXLTS U2281 ( .AN(genblk1_3__mac_biasesStored[0]), .B(n2125), .Y(n48)
         );
  NAND2BXLTS U2282 ( .AN(genblk1_0__mac_biasesStored[0]), .B(n2124), .Y(n12)
         );
  NAND2BXLTS U2283 ( .AN(genblk1_2__mac_biasesStored[0]), .B(n2125), .Y(n36)
         );
  CLKBUFX2TS U2284 ( .A(n2133), .Y(n2126) );
  CLKBUFX2TS U2285 ( .A(n2126), .Y(n2143) );
  CLKBUFX2TS U2286 ( .A(n2126), .Y(n2144) );
  CLKBUFX2TS U2287 ( .A(n2126), .Y(n2145) );
  NAND2BXLTS U2288 ( .AN(genblk1_8__mac_biasesStored[0]), .B(n2127), .Y(n108)
         );
  NAND2BXLTS U2289 ( .AN(genblk1_5__mac_biasesStored[0]), .B(n2128), .Y(n72)
         );
  NAND2BXLTS U2290 ( .AN(genblk1_4__mac_biasesStored[0]), .B(n2128), .Y(n60)
         );
  CLKBUFX2TS U2291 ( .A(n2129), .Y(n2136) );
  CLKBUFX2TS U2292 ( .A(n2129), .Y(n2138) );
endmodule

