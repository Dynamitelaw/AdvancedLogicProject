
module Layer2WeightStorage ( writeEnable, NodeSelect, writeIn, readOut );
  input [2:0] NodeSelect;
  input [59:0] writeIn;
  output [59:0] readOut;
  input writeEnable;
  wire   n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
  wire   [479:0] readOutBus;

  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_40_ ( .G(n934), .D(n847), .Q(
        readOutBus[160]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_41_ ( .G(n934), .D(n849), .Q(
        readOutBus[161]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_42_ ( .G(n934), .D(n851), .Q(
        readOutBus[162]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_43_ ( .G(n934), .D(n853), .Q(
        readOutBus[163]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_44_ ( .G(n933), .D(n855), .Q(
        readOutBus[164]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_45_ ( .G(n933), .D(n857), .Q(
        readOutBus[165]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_46_ ( .G(n933), .D(n859), .Q(
        readOutBus[166]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_47_ ( .G(n933), .D(n861), .Q(
        readOutBus[167]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_48_ ( .G(n932), .D(n863), .Q(
        readOutBus[168]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_49_ ( .G(n932), .D(n865), .Q(
        readOutBus[169]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_50_ ( .G(n932), .D(n867), .Q(
        readOutBus[170]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_51_ ( .G(n932), .D(n869), .Q(
        readOutBus[171]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_52_ ( .G(n931), .D(n871), .Q(
        readOutBus[172]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_53_ ( .G(n931), .D(n873), .Q(
        readOutBus[173]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_54_ ( .G(n931), .D(n875), .Q(
        readOutBus[174]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_55_ ( .G(n931), .D(n877), .Q(
        readOutBus[175]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_56_ ( .G(n930), .D(n879), .Q(
        readOutBus[176]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_57_ ( .G(n930), .D(n881), .Q(
        readOutBus[177]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_58_ ( .G(n930), .D(n883), .Q(
        readOutBus[178]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_59_ ( .G(n930), .D(n885), .Q(
        readOutBus[179]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_36_ ( .G(n948), .D(n839), .Q(
        readOutBus[216]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_37_ ( .G(n948), .D(n841), .Q(
        readOutBus[217]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_38_ ( .G(n948), .D(n843), .Q(
        readOutBus[218]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_39_ ( .G(n948), .D(n845), .Q(
        readOutBus[219]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_44_ ( .G(n354), .D(n855), .Q(
        readOutBus[224]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_45_ ( .G(n355), .D(n857), .Q(
        readOutBus[225]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_46_ ( .G(n327), .D(n859), .Q(
        readOutBus[226]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_47_ ( .G(n327), .D(n861), .Q(
        readOutBus[227]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_40_ ( .G(n989), .D(n847), .Q(
        readOutBus[400]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_41_ ( .G(n989), .D(n849), .Q(
        readOutBus[401]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_42_ ( .G(n989), .D(n851), .Q(
        readOutBus[402]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_43_ ( .G(n989), .D(n853), .Q(
        readOutBus[403]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_44_ ( .G(n988), .D(n855), .Q(
        readOutBus[404]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_45_ ( .G(n988), .D(n857), .Q(
        readOutBus[405]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_46_ ( .G(n988), .D(n859), .Q(
        readOutBus[406]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_47_ ( .G(n988), .D(n861), .Q(
        readOutBus[407]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_48_ ( .G(n987), .D(n863), .Q(
        readOutBus[408]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_49_ ( .G(n987), .D(n865), .Q(
        readOutBus[409]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_50_ ( .G(n987), .D(n867), .Q(
        readOutBus[410]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_51_ ( .G(n987), .D(n869), .Q(
        readOutBus[411]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_52_ ( .G(n986), .D(n871), .Q(
        readOutBus[412]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_53_ ( .G(n986), .D(n873), .Q(
        readOutBus[413]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_54_ ( .G(n986), .D(n875), .Q(
        readOutBus[414]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_55_ ( .G(n986), .D(n877), .Q(
        readOutBus[415]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_56_ ( .G(n985), .D(n879), .Q(
        readOutBus[416]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_57_ ( .G(n985), .D(n881), .Q(
        readOutBus[417]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_58_ ( .G(n985), .D(n883), .Q(
        readOutBus[418]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_59_ ( .G(n985), .D(n885), .Q(
        readOutBus[419]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_36_ ( .G(n1003), .D(n839), 
        .Q(readOutBus[456]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_37_ ( .G(n1003), .D(n841), 
        .Q(readOutBus[457]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_38_ ( .G(n1003), .D(n843), 
        .Q(readOutBus[458]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_39_ ( .G(n1003), .D(n845), 
        .Q(readOutBus[459]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_44_ ( .G(n358), .D(n855), .Q(
        readOutBus[464]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_45_ ( .G(n359), .D(n857), .Q(
        readOutBus[465]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_46_ ( .G(n321), .D(n859), .Q(
        readOutBus[466]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_47_ ( .G(n321), .D(n861), .Q(
        readOutBus[467]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_0_ ( .G(n943), .D(n767), .Q(
        readOutBus[120]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_1_ ( .G(n943), .D(n769), .Q(
        readOutBus[121]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_2_ ( .G(n943), .D(n771), .Q(
        readOutBus[122]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_3_ ( .G(n943), .D(n773), .Q(
        readOutBus[123]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_8_ ( .G(n942), .D(n783), .Q(
        readOutBus[128]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_9_ ( .G(n942), .D(n785), .Q(
        readOutBus[129]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_10_ ( .G(n942), .D(n787), .Q(
        readOutBus[130]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_11_ ( .G(n942), .D(n789), .Q(
        readOutBus[131]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_0_ ( .G(n956), .D(n767), .Q(
        readOutBus[180]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_1_ ( .G(n956), .D(n769), .Q(
        readOutBus[181]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_2_ ( .G(n956), .D(n771), .Q(
        readOutBus[182]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_3_ ( .G(n956), .D(n773), .Q(
        readOutBus[183]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_8_ ( .G(n955), .D(n783), .Q(
        readOutBus[188]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_9_ ( .G(n955), .D(n785), .Q(
        readOutBus[189]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_10_ ( .G(n955), .D(n787), .Q(
        readOutBus[190]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_11_ ( .G(n955), .D(n789), .Q(
        readOutBus[191]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_0_ ( .G(n998), .D(n767), .Q(
        readOutBus[360]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_1_ ( .G(n998), .D(n769), .Q(
        readOutBus[361]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_2_ ( .G(n998), .D(n771), .Q(
        readOutBus[362]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_3_ ( .G(n998), .D(n773), .Q(
        readOutBus[363]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_8_ ( .G(n997), .D(n783), .Q(
        readOutBus[368]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_9_ ( .G(n997), .D(n785), .Q(
        readOutBus[369]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_10_ ( .G(n997), .D(n787), .Q(
        readOutBus[370]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_11_ ( .G(n997), .D(n789), .Q(
        readOutBus[371]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_0_ ( .G(n1011), .D(n767), .Q(
        readOutBus[420]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_1_ ( .G(n1011), .D(n769), .Q(
        readOutBus[421]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_2_ ( .G(n1011), .D(n771), .Q(
        readOutBus[422]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_3_ ( .G(n1011), .D(n773), .Q(
        readOutBus[423]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_8_ ( .G(n1010), .D(n783), .Q(
        readOutBus[428]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_9_ ( .G(n1010), .D(n785), .Q(
        readOutBus[429]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_10_ ( .G(n1010), .D(n787), 
        .Q(readOutBus[430]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_11_ ( .G(n1010), .D(n789), 
        .Q(readOutBus[431]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_12_ ( .G(n941), .D(n791), .Q(
        readOutBus[132]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_13_ ( .G(n941), .D(n793), .Q(
        readOutBus[133]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_14_ ( .G(n941), .D(n795), .Q(
        readOutBus[134]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_15_ ( .G(n941), .D(n797), .Q(
        readOutBus[135]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_16_ ( .G(n940), .D(n799), .Q(
        readOutBus[136]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_17_ ( .G(n940), .D(n801), .Q(
        readOutBus[137]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_18_ ( .G(n940), .D(n803), .Q(
        readOutBus[138]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_19_ ( .G(n940), .D(n805), .Q(
        readOutBus[139]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_20_ ( .G(n939), .D(n807), .Q(
        readOutBus[140]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_21_ ( .G(n939), .D(n809), .Q(
        readOutBus[141]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_22_ ( .G(n939), .D(n811), .Q(
        readOutBus[142]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_23_ ( .G(n939), .D(n813), .Q(
        readOutBus[143]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_24_ ( .G(n938), .D(n815), .Q(
        readOutBus[144]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_25_ ( .G(n938), .D(n817), .Q(
        readOutBus[145]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_26_ ( .G(n938), .D(n819), .Q(
        readOutBus[146]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_27_ ( .G(n938), .D(n821), .Q(
        readOutBus[147]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_28_ ( .G(n937), .D(n823), .Q(
        readOutBus[148]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_29_ ( .G(n937), .D(n825), .Q(
        readOutBus[149]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_30_ ( .G(n937), .D(n827), .Q(
        readOutBus[150]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_31_ ( .G(n937), .D(n829), .Q(
        readOutBus[151]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_32_ ( .G(n936), .D(n831), .Q(
        readOutBus[152]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_33_ ( .G(n936), .D(n833), .Q(
        readOutBus[153]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_34_ ( .G(n936), .D(n835), .Q(
        readOutBus[154]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_35_ ( .G(n936), .D(n837), .Q(
        readOutBus[155]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_36_ ( .G(n935), .D(n839), .Q(
        readOutBus[156]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_37_ ( .G(n935), .D(n841), .Q(
        readOutBus[157]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_38_ ( .G(n935), .D(n843), .Q(
        readOutBus[158]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_39_ ( .G(n935), .D(n845), .Q(
        readOutBus[159]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_12_ ( .G(n954), .D(n791), .Q(
        readOutBus[192]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_13_ ( .G(n954), .D(n793), .Q(
        readOutBus[193]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_14_ ( .G(n954), .D(n795), .Q(
        readOutBus[194]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_15_ ( .G(n954), .D(n797), .Q(
        readOutBus[195]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_16_ ( .G(n953), .D(n799), .Q(
        readOutBus[196]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_17_ ( .G(n953), .D(n801), .Q(
        readOutBus[197]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_18_ ( .G(n953), .D(n803), .Q(
        readOutBus[198]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_19_ ( .G(n953), .D(n805), .Q(
        readOutBus[199]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_20_ ( .G(n952), .D(n807), .Q(
        readOutBus[200]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_21_ ( .G(n952), .D(n809), .Q(
        readOutBus[201]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_22_ ( .G(n952), .D(n811), .Q(
        readOutBus[202]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_23_ ( .G(n952), .D(n813), .Q(
        readOutBus[203]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_24_ ( .G(n951), .D(n815), .Q(
        readOutBus[204]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_25_ ( .G(n951), .D(n817), .Q(
        readOutBus[205]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_26_ ( .G(n951), .D(n819), .Q(
        readOutBus[206]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_27_ ( .G(n951), .D(n821), .Q(
        readOutBus[207]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_28_ ( .G(n950), .D(n823), .Q(
        readOutBus[208]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_29_ ( .G(n950), .D(n825), .Q(
        readOutBus[209]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_30_ ( .G(n950), .D(n827), .Q(
        readOutBus[210]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_31_ ( .G(n950), .D(n829), .Q(
        readOutBus[211]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_32_ ( .G(n949), .D(n831), .Q(
        readOutBus[212]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_33_ ( .G(n949), .D(n833), .Q(
        readOutBus[213]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_34_ ( .G(n949), .D(n835), .Q(
        readOutBus[214]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_35_ ( .G(n949), .D(n837), .Q(
        readOutBus[215]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_40_ ( .G(n947), .D(n847), .Q(
        readOutBus[220]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_41_ ( .G(n947), .D(n849), .Q(
        readOutBus[221]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_42_ ( .G(n947), .D(n851), .Q(
        readOutBus[222]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_43_ ( .G(n947), .D(n853), .Q(
        readOutBus[223]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_48_ ( .G(n946), .D(n863), .Q(
        readOutBus[228]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_49_ ( .G(n946), .D(n865), .Q(
        readOutBus[229]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_50_ ( .G(n946), .D(n867), .Q(
        readOutBus[230]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_51_ ( .G(n946), .D(n869), .Q(
        readOutBus[231]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_52_ ( .G(n945), .D(n871), .Q(
        readOutBus[232]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_53_ ( .G(n945), .D(n873), .Q(
        readOutBus[233]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_54_ ( .G(n945), .D(n875), .Q(
        readOutBus[234]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_55_ ( .G(n945), .D(n877), .Q(
        readOutBus[235]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_56_ ( .G(n944), .D(n879), .Q(
        readOutBus[236]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_57_ ( .G(n944), .D(n881), .Q(
        readOutBus[237]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_58_ ( .G(n944), .D(n883), .Q(
        readOutBus[238]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_59_ ( .G(n944), .D(n885), .Q(
        readOutBus[239]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_12_ ( .G(n996), .D(n791), .Q(
        readOutBus[372]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_13_ ( .G(n996), .D(n793), .Q(
        readOutBus[373]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_14_ ( .G(n996), .D(n795), .Q(
        readOutBus[374]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_15_ ( .G(n996), .D(n797), .Q(
        readOutBus[375]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_16_ ( .G(n995), .D(n799), .Q(
        readOutBus[376]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_17_ ( .G(n995), .D(n801), .Q(
        readOutBus[377]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_18_ ( .G(n995), .D(n803), .Q(
        readOutBus[378]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_19_ ( .G(n995), .D(n805), .Q(
        readOutBus[379]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_20_ ( .G(n994), .D(n807), .Q(
        readOutBus[380]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_21_ ( .G(n994), .D(n809), .Q(
        readOutBus[381]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_22_ ( .G(n994), .D(n811), .Q(
        readOutBus[382]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_23_ ( .G(n994), .D(n813), .Q(
        readOutBus[383]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_24_ ( .G(n993), .D(n815), .Q(
        readOutBus[384]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_25_ ( .G(n993), .D(n817), .Q(
        readOutBus[385]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_26_ ( .G(n993), .D(n819), .Q(
        readOutBus[386]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_27_ ( .G(n993), .D(n821), .Q(
        readOutBus[387]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_28_ ( .G(n992), .D(n823), .Q(
        readOutBus[388]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_29_ ( .G(n992), .D(n825), .Q(
        readOutBus[389]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_30_ ( .G(n992), .D(n827), .Q(
        readOutBus[390]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_31_ ( .G(n992), .D(n829), .Q(
        readOutBus[391]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_32_ ( .G(n991), .D(n831), .Q(
        readOutBus[392]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_33_ ( .G(n991), .D(n833), .Q(
        readOutBus[393]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_34_ ( .G(n991), .D(n835), .Q(
        readOutBus[394]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_35_ ( .G(n991), .D(n837), .Q(
        readOutBus[395]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_36_ ( .G(n990), .D(n839), .Q(
        readOutBus[396]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_37_ ( .G(n990), .D(n841), .Q(
        readOutBus[397]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_38_ ( .G(n990), .D(n843), .Q(
        readOutBus[398]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_39_ ( .G(n990), .D(n845), .Q(
        readOutBus[399]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_12_ ( .G(n1009), .D(n791), 
        .Q(readOutBus[432]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_13_ ( .G(n1009), .D(n793), 
        .Q(readOutBus[433]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_14_ ( .G(n1009), .D(n795), 
        .Q(readOutBus[434]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_15_ ( .G(n1009), .D(n797), 
        .Q(readOutBus[435]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_16_ ( .G(n1008), .D(n799), 
        .Q(readOutBus[436]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_17_ ( .G(n1008), .D(n801), 
        .Q(readOutBus[437]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_18_ ( .G(n1008), .D(n803), 
        .Q(readOutBus[438]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_19_ ( .G(n1008), .D(n805), 
        .Q(readOutBus[439]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_20_ ( .G(n1007), .D(n807), 
        .Q(readOutBus[440]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_21_ ( .G(n1007), .D(n809), 
        .Q(readOutBus[441]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_22_ ( .G(n1007), .D(n811), 
        .Q(readOutBus[442]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_23_ ( .G(n1007), .D(n813), 
        .Q(readOutBus[443]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_24_ ( .G(n1006), .D(n815), 
        .Q(readOutBus[444]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_25_ ( .G(n1006), .D(n817), 
        .Q(readOutBus[445]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_26_ ( .G(n1006), .D(n819), 
        .Q(readOutBus[446]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_27_ ( .G(n1006), .D(n821), 
        .Q(readOutBus[447]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_28_ ( .G(n1005), .D(n823), 
        .Q(readOutBus[448]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_29_ ( .G(n1005), .D(n825), 
        .Q(readOutBus[449]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_30_ ( .G(n1005), .D(n827), 
        .Q(readOutBus[450]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_31_ ( .G(n1005), .D(n829), 
        .Q(readOutBus[451]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_32_ ( .G(n1004), .D(n831), 
        .Q(readOutBus[452]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_33_ ( .G(n1004), .D(n833), 
        .Q(readOutBus[453]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_34_ ( .G(n1004), .D(n835), 
        .Q(readOutBus[454]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_35_ ( .G(n1004), .D(n837), 
        .Q(readOutBus[455]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_40_ ( .G(n1002), .D(n847), 
        .Q(readOutBus[460]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_41_ ( .G(n1002), .D(n849), 
        .Q(readOutBus[461]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_42_ ( .G(n1002), .D(n851), 
        .Q(readOutBus[462]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_43_ ( .G(n1002), .D(n853), 
        .Q(readOutBus[463]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_48_ ( .G(n1001), .D(n863), 
        .Q(readOutBus[468]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_49_ ( .G(n1001), .D(n865), 
        .Q(readOutBus[469]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_50_ ( .G(n1001), .D(n867), 
        .Q(readOutBus[470]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_51_ ( .G(n1001), .D(n869), 
        .Q(readOutBus[471]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_52_ ( .G(n1000), .D(n871), 
        .Q(readOutBus[472]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_53_ ( .G(n1000), .D(n873), 
        .Q(readOutBus[473]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_54_ ( .G(n1000), .D(n875), 
        .Q(readOutBus[474]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_55_ ( .G(n1000), .D(n877), 
        .Q(readOutBus[475]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_56_ ( .G(n999), .D(n879), .Q(
        readOutBus[476]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_57_ ( .G(n999), .D(n881), .Q(
        readOutBus[477]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_58_ ( .G(n999), .D(n883), .Q(
        readOutBus[478]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_59_ ( .G(n999), .D(n885), .Q(
        readOutBus[479]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_5_ ( .G(n890), .D(n777), .Q(
        readOutBus[125]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_7_ ( .G(n890), .D(n781), .Q(
        readOutBus[127]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_5_ ( .G(n898), .D(n777), .Q(
        readOutBus[365]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_7_ ( .G(n898), .D(n781), .Q(
        readOutBus[367]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_5_ ( .G(n892), .D(n777), .Q(
        readOutBus[185]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_7_ ( .G(n892), .D(n781), .Q(
        readOutBus[187]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_5_ ( .G(n900), .D(n777), .Q(
        readOutBus[425]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_7_ ( .G(n900), .D(n781), .Q(
        readOutBus[427]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_4_ ( .G(n891), .D(n775), .Q(
        readOutBus[124]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_6_ ( .G(n891), .D(n779), .Q(
        readOutBus[126]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_4_ ( .G(n893), .D(n775), .Q(
        readOutBus[184]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_6_ ( .G(n893), .D(n779), .Q(
        readOutBus[186]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_4_ ( .G(n899), .D(n775), .Q(
        readOutBus[364]) );
  TLATXLTS Generate_Node_Banks_6__NB_readOut_reg_6_ ( .G(n899), .D(n779), .Q(
        readOutBus[366]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_4_ ( .G(n901), .D(n775), .Q(
        readOutBus[424]) );
  TLATXLTS Generate_Node_Banks_7__NB_readOut_reg_6_ ( .G(n901), .D(n779), .Q(
        readOutBus[426]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_40_ ( .G(n906), .D(n846), .Q(
        readOutBus[40]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_41_ ( .G(n906), .D(n848), .Q(
        readOutBus[41]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_42_ ( .G(n906), .D(n850), .Q(
        readOutBus[42]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_43_ ( .G(n906), .D(n852), .Q(
        readOutBus[43]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_44_ ( .G(n905), .D(n854), .Q(
        readOutBus[44]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_45_ ( .G(n905), .D(n856), .Q(
        readOutBus[45]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_46_ ( .G(n905), .D(n858), .Q(
        readOutBus[46]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_47_ ( .G(n905), .D(n860), .Q(
        readOutBus[47]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_48_ ( .G(n904), .D(n862), .Q(
        readOutBus[48]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_49_ ( .G(n904), .D(n864), .Q(
        readOutBus[49]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_50_ ( .G(n904), .D(n866), .Q(
        readOutBus[50]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_51_ ( .G(n904), .D(n868), .Q(
        readOutBus[51]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_52_ ( .G(n903), .D(n870), .Q(
        readOutBus[52]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_53_ ( .G(n903), .D(n872), .Q(
        readOutBus[53]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_54_ ( .G(n903), .D(n874), .Q(
        readOutBus[54]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_55_ ( .G(n903), .D(n876), .Q(
        readOutBus[55]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_56_ ( .G(n902), .D(n878), .Q(
        readOutBus[56]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_57_ ( .G(n902), .D(n880), .Q(
        readOutBus[57]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_58_ ( .G(n902), .D(n882), .Q(
        readOutBus[58]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_59_ ( .G(n902), .D(n884), .Q(
        readOutBus[59]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_40_ ( .G(n920), .D(n846), .Q(
        readOutBus[100]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_41_ ( .G(n920), .D(n848), .Q(
        readOutBus[101]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_42_ ( .G(n920), .D(n850), .Q(
        readOutBus[102]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_43_ ( .G(n920), .D(n852), .Q(
        readOutBus[103]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_44_ ( .G(n919), .D(n854), .Q(
        readOutBus[104]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_45_ ( .G(n919), .D(n856), .Q(
        readOutBus[105]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_46_ ( .G(n919), .D(n858), .Q(
        readOutBus[106]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_47_ ( .G(n919), .D(n860), .Q(
        readOutBus[107]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_48_ ( .G(n918), .D(n862), .Q(
        readOutBus[108]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_49_ ( .G(n918), .D(n864), .Q(
        readOutBus[109]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_50_ ( .G(n918), .D(n866), .Q(
        readOutBus[110]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_51_ ( .G(n918), .D(n868), .Q(
        readOutBus[111]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_52_ ( .G(n917), .D(n870), .Q(
        readOutBus[112]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_53_ ( .G(n917), .D(n872), .Q(
        readOutBus[113]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_54_ ( .G(n917), .D(n874), .Q(
        readOutBus[114]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_55_ ( .G(n917), .D(n876), .Q(
        readOutBus[115]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_56_ ( .G(n916), .D(n878), .Q(
        readOutBus[116]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_57_ ( .G(n916), .D(n880), .Q(
        readOutBus[117]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_58_ ( .G(n916), .D(n882), .Q(
        readOutBus[118]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_59_ ( .G(n916), .D(n884), .Q(
        readOutBus[119]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_40_ ( .G(n961), .D(n846), .Q(
        readOutBus[280]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_41_ ( .G(n961), .D(n848), .Q(
        readOutBus[281]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_42_ ( .G(n961), .D(n850), .Q(
        readOutBus[282]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_43_ ( .G(n961), .D(n852), .Q(
        readOutBus[283]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_44_ ( .G(n960), .D(n854), .Q(
        readOutBus[284]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_45_ ( .G(n960), .D(n856), .Q(
        readOutBus[285]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_46_ ( .G(n960), .D(n858), .Q(
        readOutBus[286]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_47_ ( .G(n960), .D(n860), .Q(
        readOutBus[287]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_48_ ( .G(n959), .D(n862), .Q(
        readOutBus[288]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_49_ ( .G(n959), .D(n864), .Q(
        readOutBus[289]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_50_ ( .G(n959), .D(n866), .Q(
        readOutBus[290]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_51_ ( .G(n959), .D(n868), .Q(
        readOutBus[291]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_52_ ( .G(n958), .D(n870), .Q(
        readOutBus[292]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_53_ ( .G(n958), .D(n872), .Q(
        readOutBus[293]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_54_ ( .G(n958), .D(n874), .Q(
        readOutBus[294]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_55_ ( .G(n958), .D(n876), .Q(
        readOutBus[295]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_56_ ( .G(n957), .D(n878), .Q(
        readOutBus[296]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_57_ ( .G(n957), .D(n880), .Q(
        readOutBus[297]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_58_ ( .G(n957), .D(n882), .Q(
        readOutBus[298]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_59_ ( .G(n957), .D(n884), .Q(
        readOutBus[299]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_40_ ( .G(n975), .D(n846), .Q(
        readOutBus[340]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_41_ ( .G(n975), .D(n848), .Q(
        readOutBus[341]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_42_ ( .G(n975), .D(n850), .Q(
        readOutBus[342]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_43_ ( .G(n975), .D(n852), .Q(
        readOutBus[343]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_44_ ( .G(n974), .D(n854), .Q(
        readOutBus[344]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_45_ ( .G(n974), .D(n856), .Q(
        readOutBus[345]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_46_ ( .G(n974), .D(n858), .Q(
        readOutBus[346]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_47_ ( .G(n974), .D(n860), .Q(
        readOutBus[347]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_48_ ( .G(n973), .D(n862), .Q(
        readOutBus[348]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_49_ ( .G(n973), .D(n864), .Q(
        readOutBus[349]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_50_ ( .G(n973), .D(n866), .Q(
        readOutBus[350]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_51_ ( .G(n973), .D(n868), .Q(
        readOutBus[351]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_52_ ( .G(n972), .D(n870), .Q(
        readOutBus[352]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_53_ ( .G(n972), .D(n872), .Q(
        readOutBus[353]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_54_ ( .G(n972), .D(n874), .Q(
        readOutBus[354]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_55_ ( .G(n972), .D(n876), .Q(
        readOutBus[355]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_56_ ( .G(n971), .D(n878), .Q(
        readOutBus[356]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_57_ ( .G(n971), .D(n880), .Q(
        readOutBus[357]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_58_ ( .G(n971), .D(n882), .Q(
        readOutBus[358]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_59_ ( .G(n971), .D(n884), .Q(
        readOutBus[359]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_24_ ( .G(n910), .D(n814), .Q(
        readOutBus[24]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_25_ ( .G(n910), .D(n816), .Q(
        readOutBus[25]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_26_ ( .G(n910), .D(n818), .Q(
        readOutBus[26]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_27_ ( .G(n910), .D(n820), .Q(
        readOutBus[27]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_28_ ( .G(n909), .D(n822), .Q(
        readOutBus[28]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_29_ ( .G(n909), .D(n824), .Q(
        readOutBus[29]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_30_ ( .G(n909), .D(n826), .Q(
        readOutBus[30]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_31_ ( .G(n909), .D(n828), .Q(
        readOutBus[31]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_32_ ( .G(n908), .D(n830), .Q(
        readOutBus[32]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_33_ ( .G(n908), .D(n832), .Q(
        readOutBus[33]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_34_ ( .G(n908), .D(n834), .Q(
        readOutBus[34]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_35_ ( .G(n908), .D(n836), .Q(
        readOutBus[35]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_36_ ( .G(n907), .D(n838), .Q(
        readOutBus[36]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_37_ ( .G(n907), .D(n840), .Q(
        readOutBus[37]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_38_ ( .G(n907), .D(n842), .Q(
        readOutBus[38]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_39_ ( .G(n907), .D(n844), .Q(
        readOutBus[39]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_24_ ( .G(n924), .D(n814), .Q(
        readOutBus[84]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_25_ ( .G(n924), .D(n816), .Q(
        readOutBus[85]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_26_ ( .G(n924), .D(n818), .Q(
        readOutBus[86]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_27_ ( .G(n924), .D(n820), .Q(
        readOutBus[87]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_28_ ( .G(n923), .D(n822), .Q(
        readOutBus[88]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_29_ ( .G(n923), .D(n824), .Q(
        readOutBus[89]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_30_ ( .G(n923), .D(n826), .Q(
        readOutBus[90]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_31_ ( .G(n923), .D(n828), .Q(
        readOutBus[91]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_32_ ( .G(n922), .D(n830), .Q(
        readOutBus[92]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_33_ ( .G(n922), .D(n832), .Q(
        readOutBus[93]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_34_ ( .G(n922), .D(n834), .Q(
        readOutBus[94]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_35_ ( .G(n922), .D(n836), .Q(
        readOutBus[95]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_36_ ( .G(n921), .D(n838), .Q(
        readOutBus[96]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_37_ ( .G(n921), .D(n840), .Q(
        readOutBus[97]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_38_ ( .G(n921), .D(n842), .Q(
        readOutBus[98]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_39_ ( .G(n921), .D(n844), .Q(
        readOutBus[99]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_24_ ( .G(n965), .D(n814), .Q(
        readOutBus[264]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_25_ ( .G(n965), .D(n816), .Q(
        readOutBus[265]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_26_ ( .G(n965), .D(n818), .Q(
        readOutBus[266]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_27_ ( .G(n965), .D(n820), .Q(
        readOutBus[267]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_28_ ( .G(n964), .D(n822), .Q(
        readOutBus[268]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_29_ ( .G(n964), .D(n824), .Q(
        readOutBus[269]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_30_ ( .G(n964), .D(n826), .Q(
        readOutBus[270]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_31_ ( .G(n964), .D(n828), .Q(
        readOutBus[271]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_32_ ( .G(n963), .D(n830), .Q(
        readOutBus[272]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_33_ ( .G(n963), .D(n832), .Q(
        readOutBus[273]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_34_ ( .G(n963), .D(n834), .Q(
        readOutBus[274]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_35_ ( .G(n963), .D(n836), .Q(
        readOutBus[275]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_36_ ( .G(n962), .D(n838), .Q(
        readOutBus[276]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_37_ ( .G(n962), .D(n840), .Q(
        readOutBus[277]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_38_ ( .G(n962), .D(n842), .Q(
        readOutBus[278]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_39_ ( .G(n962), .D(n844), .Q(
        readOutBus[279]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_24_ ( .G(n979), .D(n814), .Q(
        readOutBus[324]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_25_ ( .G(n979), .D(n816), .Q(
        readOutBus[325]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_26_ ( .G(n979), .D(n818), .Q(
        readOutBus[326]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_27_ ( .G(n979), .D(n820), .Q(
        readOutBus[327]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_28_ ( .G(n978), .D(n822), .Q(
        readOutBus[328]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_29_ ( .G(n978), .D(n824), .Q(
        readOutBus[329]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_30_ ( .G(n978), .D(n826), .Q(
        readOutBus[330]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_31_ ( .G(n978), .D(n828), .Q(
        readOutBus[331]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_32_ ( .G(n977), .D(n830), .Q(
        readOutBus[332]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_33_ ( .G(n977), .D(n832), .Q(
        readOutBus[333]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_34_ ( .G(n977), .D(n834), .Q(
        readOutBus[334]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_35_ ( .G(n977), .D(n836), .Q(
        readOutBus[335]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_36_ ( .G(n976), .D(n838), .Q(
        readOutBus[336]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_37_ ( .G(n976), .D(n840), .Q(
        readOutBus[337]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_38_ ( .G(n976), .D(n842), .Q(
        readOutBus[338]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_39_ ( .G(n976), .D(n844), .Q(
        readOutBus[339]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_0_ ( .G(n915), .D(n766), .Q(
        readOutBus[0]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_1_ ( .G(n915), .D(n768), .Q(
        readOutBus[1]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_2_ ( .G(n915), .D(n770), .Q(
        readOutBus[2]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_3_ ( .G(n915), .D(n772), .Q(
        readOutBus[3]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_8_ ( .G(n914), .D(n782), .Q(
        readOutBus[8]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_9_ ( .G(n914), .D(n784), .Q(
        readOutBus[9]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_10_ ( .G(n914), .D(n786), .Q(
        readOutBus[10]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_11_ ( .G(n914), .D(n788), .Q(
        readOutBus[11]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_0_ ( .G(n929), .D(n766), .Q(
        readOutBus[60]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_1_ ( .G(n929), .D(n768), .Q(
        readOutBus[61]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_2_ ( .G(n929), .D(n770), .Q(
        readOutBus[62]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_3_ ( .G(n929), .D(n772), .Q(
        readOutBus[63]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_8_ ( .G(n928), .D(n782), .Q(
        readOutBus[68]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_9_ ( .G(n928), .D(n784), .Q(
        readOutBus[69]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_10_ ( .G(n928), .D(n786), .Q(
        readOutBus[70]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_11_ ( .G(n928), .D(n788), .Q(
        readOutBus[71]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_0_ ( .G(n970), .D(n766), .Q(
        readOutBus[240]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_1_ ( .G(n970), .D(n768), .Q(
        readOutBus[241]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_2_ ( .G(n970), .D(n770), .Q(
        readOutBus[242]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_3_ ( .G(n970), .D(n772), .Q(
        readOutBus[243]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_8_ ( .G(n969), .D(n782), .Q(
        readOutBus[248]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_9_ ( .G(n969), .D(n784), .Q(
        readOutBus[249]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_10_ ( .G(n969), .D(n786), .Q(
        readOutBus[250]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_11_ ( .G(n969), .D(n788), .Q(
        readOutBus[251]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_0_ ( .G(n984), .D(n766), .Q(
        readOutBus[300]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_1_ ( .G(n984), .D(n768), .Q(
        readOutBus[301]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_2_ ( .G(n984), .D(n770), .Q(
        readOutBus[302]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_3_ ( .G(n984), .D(n772), .Q(
        readOutBus[303]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_8_ ( .G(n983), .D(n782), .Q(
        readOutBus[308]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_9_ ( .G(n983), .D(n784), .Q(
        readOutBus[309]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_10_ ( .G(n983), .D(n786), .Q(
        readOutBus[310]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_11_ ( .G(n983), .D(n788), .Q(
        readOutBus[311]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_5_ ( .G(n886), .D(n776), .Q(
        readOutBus[5]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_7_ ( .G(n886), .D(n780), .Q(
        readOutBus[7]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_5_ ( .G(n888), .D(n776), .Q(
        readOutBus[65]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_7_ ( .G(n888), .D(n780), .Q(
        readOutBus[67]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_5_ ( .G(n894), .D(n776), .Q(
        readOutBus[245]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_7_ ( .G(n894), .D(n780), .Q(
        readOutBus[247]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_5_ ( .G(n896), .D(n776), .Q(
        readOutBus[305]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_7_ ( .G(n896), .D(n780), .Q(
        readOutBus[307]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_12_ ( .G(n913), .D(n790), .Q(
        readOutBus[12]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_13_ ( .G(n913), .D(n792), .Q(
        readOutBus[13]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_14_ ( .G(n913), .D(n794), .Q(
        readOutBus[14]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_15_ ( .G(n913), .D(n796), .Q(
        readOutBus[15]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_16_ ( .G(n912), .D(n798), .Q(
        readOutBus[16]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_17_ ( .G(n912), .D(n800), .Q(
        readOutBus[17]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_18_ ( .G(n912), .D(n802), .Q(
        readOutBus[18]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_19_ ( .G(n912), .D(n804), .Q(
        readOutBus[19]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_20_ ( .G(n911), .D(n806), .Q(
        readOutBus[20]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_21_ ( .G(n911), .D(n808), .Q(
        readOutBus[21]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_22_ ( .G(n911), .D(n810), .Q(
        readOutBus[22]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_23_ ( .G(n911), .D(n812), .Q(
        readOutBus[23]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_12_ ( .G(n927), .D(n790), .Q(
        readOutBus[72]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_13_ ( .G(n927), .D(n792), .Q(
        readOutBus[73]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_14_ ( .G(n927), .D(n794), .Q(
        readOutBus[74]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_15_ ( .G(n927), .D(n796), .Q(
        readOutBus[75]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_16_ ( .G(n926), .D(n798), .Q(
        readOutBus[76]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_17_ ( .G(n926), .D(n800), .Q(
        readOutBus[77]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_18_ ( .G(n926), .D(n802), .Q(
        readOutBus[78]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_19_ ( .G(n926), .D(n804), .Q(
        readOutBus[79]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_20_ ( .G(n925), .D(n806), .Q(
        readOutBus[80]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_21_ ( .G(n925), .D(n808), .Q(
        readOutBus[81]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_22_ ( .G(n925), .D(n810), .Q(
        readOutBus[82]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_23_ ( .G(n925), .D(n812), .Q(
        readOutBus[83]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_12_ ( .G(n968), .D(n790), .Q(
        readOutBus[252]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_13_ ( .G(n968), .D(n792), .Q(
        readOutBus[253]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_14_ ( .G(n968), .D(n794), .Q(
        readOutBus[254]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_15_ ( .G(n968), .D(n796), .Q(
        readOutBus[255]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_16_ ( .G(n967), .D(n798), .Q(
        readOutBus[256]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_17_ ( .G(n967), .D(n800), .Q(
        readOutBus[257]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_18_ ( .G(n967), .D(n802), .Q(
        readOutBus[258]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_19_ ( .G(n967), .D(n804), .Q(
        readOutBus[259]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_20_ ( .G(n966), .D(n806), .Q(
        readOutBus[260]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_21_ ( .G(n966), .D(n808), .Q(
        readOutBus[261]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_22_ ( .G(n966), .D(n810), .Q(
        readOutBus[262]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_23_ ( .G(n966), .D(n812), .Q(
        readOutBus[263]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_12_ ( .G(n982), .D(n790), .Q(
        readOutBus[312]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_13_ ( .G(n982), .D(n792), .Q(
        readOutBus[313]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_14_ ( .G(n982), .D(n794), .Q(
        readOutBus[314]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_15_ ( .G(n982), .D(n796), .Q(
        readOutBus[315]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_16_ ( .G(n981), .D(n798), .Q(
        readOutBus[316]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_17_ ( .G(n981), .D(n800), .Q(
        readOutBus[317]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_18_ ( .G(n981), .D(n802), .Q(
        readOutBus[318]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_19_ ( .G(n981), .D(n804), .Q(
        readOutBus[319]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_20_ ( .G(n980), .D(n806), .Q(
        readOutBus[320]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_21_ ( .G(n980), .D(n808), .Q(
        readOutBus[321]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_22_ ( .G(n980), .D(n810), .Q(
        readOutBus[322]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_23_ ( .G(n980), .D(n812), .Q(
        readOutBus[323]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_4_ ( .G(n887), .D(n774), .Q(
        readOutBus[4]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_6_ ( .G(n887), .D(n778), .Q(
        readOutBus[6]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_4_ ( .G(n889), .D(n774), .Q(
        readOutBus[64]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_6_ ( .G(n889), .D(n778), .Q(
        readOutBus[66]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_4_ ( .G(n895), .D(n774), .Q(
        readOutBus[244]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_6_ ( .G(n895), .D(n778), .Q(
        readOutBus[246]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_4_ ( .G(n897), .D(n774), .Q(
        readOutBus[304]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_6_ ( .G(n897), .D(n778), .Q(
        readOutBus[306]) );
  INVX2TS U326 ( .A(n333), .Y(n324) );
  INVX2TS U327 ( .A(n339), .Y(n332) );
  INVX2TS U328 ( .A(n320), .Y(n337) );
  INVX2TS U329 ( .A(writeIn[0]), .Y(n256) );
  INVX2TS U330 ( .A(n256), .Y(n766) );
  INVX2TS U331 ( .A(n256), .Y(n767) );
  INVX2TS U332 ( .A(writeIn[1]), .Y(n257) );
  INVX2TS U333 ( .A(n257), .Y(n768) );
  INVX2TS U334 ( .A(n257), .Y(n769) );
  INVX2TS U335 ( .A(writeIn[2]), .Y(n258) );
  INVX2TS U336 ( .A(n258), .Y(n770) );
  INVX2TS U337 ( .A(n258), .Y(n771) );
  INVX2TS U338 ( .A(writeIn[3]), .Y(n259) );
  INVX2TS U339 ( .A(n259), .Y(n772) );
  INVX2TS U340 ( .A(n259), .Y(n773) );
  INVX2TS U341 ( .A(writeIn[4]), .Y(n260) );
  INVX2TS U342 ( .A(n260), .Y(n774) );
  INVX2TS U343 ( .A(n260), .Y(n775) );
  INVX2TS U344 ( .A(writeIn[5]), .Y(n261) );
  INVX2TS U345 ( .A(n261), .Y(n776) );
  INVX2TS U346 ( .A(n261), .Y(n777) );
  INVX2TS U347 ( .A(writeIn[6]), .Y(n262) );
  INVX2TS U348 ( .A(n262), .Y(n778) );
  INVX2TS U349 ( .A(n262), .Y(n779) );
  INVX2TS U350 ( .A(writeIn[7]), .Y(n263) );
  INVX2TS U351 ( .A(n263), .Y(n780) );
  INVX2TS U352 ( .A(n263), .Y(n781) );
  INVX2TS U353 ( .A(writeIn[8]), .Y(n264) );
  INVX2TS U354 ( .A(n264), .Y(n782) );
  INVX2TS U355 ( .A(n264), .Y(n783) );
  INVX2TS U356 ( .A(writeIn[9]), .Y(n265) );
  INVX2TS U357 ( .A(n265), .Y(n784) );
  INVX2TS U358 ( .A(n265), .Y(n785) );
  INVX2TS U359 ( .A(writeIn[10]), .Y(n266) );
  INVX2TS U360 ( .A(n266), .Y(n786) );
  INVX2TS U361 ( .A(n266), .Y(n787) );
  INVX2TS U362 ( .A(writeIn[11]), .Y(n267) );
  INVX2TS U363 ( .A(n267), .Y(n788) );
  INVX2TS U364 ( .A(n267), .Y(n789) );
  INVX2TS U365 ( .A(writeIn[12]), .Y(n268) );
  INVX2TS U366 ( .A(n268), .Y(n790) );
  INVX2TS U367 ( .A(n268), .Y(n791) );
  INVX2TS U368 ( .A(writeIn[13]), .Y(n269) );
  INVX2TS U369 ( .A(n269), .Y(n792) );
  INVX2TS U370 ( .A(n269), .Y(n793) );
  INVX2TS U371 ( .A(writeIn[14]), .Y(n270) );
  INVX2TS U372 ( .A(n270), .Y(n794) );
  INVX2TS U373 ( .A(n270), .Y(n795) );
  INVX2TS U374 ( .A(writeIn[15]), .Y(n271) );
  INVX2TS U375 ( .A(n271), .Y(n796) );
  INVX2TS U376 ( .A(n271), .Y(n797) );
  INVX2TS U377 ( .A(writeIn[16]), .Y(n272) );
  INVX2TS U378 ( .A(n272), .Y(n798) );
  INVX2TS U379 ( .A(n272), .Y(n799) );
  INVX2TS U380 ( .A(writeIn[17]), .Y(n273) );
  INVX2TS U381 ( .A(n273), .Y(n800) );
  INVX2TS U382 ( .A(n273), .Y(n801) );
  INVX2TS U383 ( .A(writeIn[18]), .Y(n274) );
  INVX2TS U384 ( .A(n274), .Y(n802) );
  INVX2TS U385 ( .A(n274), .Y(n803) );
  INVX2TS U386 ( .A(writeIn[19]), .Y(n275) );
  INVX2TS U387 ( .A(n275), .Y(n804) );
  INVX2TS U388 ( .A(n275), .Y(n805) );
  INVX2TS U389 ( .A(writeIn[20]), .Y(n276) );
  INVX2TS U390 ( .A(n276), .Y(n806) );
  INVX2TS U391 ( .A(n276), .Y(n807) );
  INVX2TS U392 ( .A(writeIn[21]), .Y(n277) );
  INVX2TS U393 ( .A(n277), .Y(n808) );
  INVX2TS U394 ( .A(n277), .Y(n809) );
  INVX2TS U395 ( .A(writeIn[22]), .Y(n278) );
  INVX2TS U396 ( .A(n278), .Y(n810) );
  INVX2TS U397 ( .A(n278), .Y(n811) );
  INVX2TS U398 ( .A(writeIn[23]), .Y(n279) );
  INVX2TS U399 ( .A(n279), .Y(n812) );
  INVX2TS U400 ( .A(n279), .Y(n813) );
  INVX2TS U401 ( .A(writeIn[24]), .Y(n280) );
  INVX2TS U402 ( .A(n280), .Y(n814) );
  INVX2TS U403 ( .A(n280), .Y(n815) );
  INVX2TS U404 ( .A(writeIn[25]), .Y(n281) );
  INVX2TS U405 ( .A(n281), .Y(n816) );
  INVX2TS U406 ( .A(n281), .Y(n817) );
  INVX2TS U407 ( .A(writeIn[26]), .Y(n282) );
  INVX2TS U408 ( .A(n282), .Y(n818) );
  INVX2TS U409 ( .A(n282), .Y(n819) );
  INVX2TS U410 ( .A(writeIn[27]), .Y(n283) );
  INVX2TS U411 ( .A(n283), .Y(n820) );
  INVX2TS U412 ( .A(n283), .Y(n821) );
  INVX2TS U413 ( .A(writeIn[28]), .Y(n284) );
  INVX2TS U414 ( .A(n284), .Y(n822) );
  INVX2TS U415 ( .A(n284), .Y(n823) );
  INVX2TS U416 ( .A(writeIn[29]), .Y(n285) );
  INVX2TS U417 ( .A(n285), .Y(n824) );
  INVX2TS U418 ( .A(n285), .Y(n825) );
  INVX2TS U419 ( .A(writeIn[30]), .Y(n286) );
  INVX2TS U420 ( .A(n286), .Y(n826) );
  INVX2TS U421 ( .A(n286), .Y(n827) );
  INVX2TS U422 ( .A(writeIn[31]), .Y(n287) );
  INVX2TS U423 ( .A(n287), .Y(n828) );
  INVX2TS U424 ( .A(n287), .Y(n829) );
  INVX2TS U425 ( .A(writeIn[32]), .Y(n288) );
  INVX2TS U426 ( .A(n288), .Y(n830) );
  INVX2TS U427 ( .A(n288), .Y(n831) );
  INVX2TS U428 ( .A(writeIn[33]), .Y(n289) );
  INVX2TS U429 ( .A(n289), .Y(n832) );
  INVX2TS U430 ( .A(n289), .Y(n833) );
  INVX2TS U431 ( .A(writeIn[34]), .Y(n290) );
  INVX2TS U432 ( .A(n290), .Y(n834) );
  INVX2TS U433 ( .A(n290), .Y(n835) );
  INVX2TS U434 ( .A(writeIn[35]), .Y(n291) );
  INVX2TS U435 ( .A(n291), .Y(n836) );
  INVX2TS U436 ( .A(n291), .Y(n837) );
  INVX2TS U437 ( .A(writeIn[36]), .Y(n292) );
  INVX2TS U438 ( .A(n292), .Y(n838) );
  INVX2TS U439 ( .A(n292), .Y(n839) );
  INVX2TS U440 ( .A(writeIn[37]), .Y(n293) );
  INVX2TS U441 ( .A(n293), .Y(n840) );
  INVX2TS U442 ( .A(n293), .Y(n841) );
  INVX2TS U443 ( .A(writeIn[38]), .Y(n294) );
  INVX2TS U444 ( .A(n294), .Y(n842) );
  INVX2TS U445 ( .A(n294), .Y(n843) );
  INVX2TS U446 ( .A(writeIn[39]), .Y(n295) );
  INVX2TS U447 ( .A(n295), .Y(n844) );
  INVX2TS U448 ( .A(n295), .Y(n845) );
  INVX2TS U449 ( .A(writeIn[40]), .Y(n296) );
  INVX2TS U450 ( .A(n296), .Y(n846) );
  INVX2TS U451 ( .A(n296), .Y(n847) );
  INVX2TS U452 ( .A(writeIn[41]), .Y(n297) );
  INVX2TS U453 ( .A(n297), .Y(n848) );
  INVX2TS U454 ( .A(n297), .Y(n849) );
  INVX2TS U455 ( .A(writeIn[42]), .Y(n298) );
  INVX2TS U456 ( .A(n298), .Y(n850) );
  INVX2TS U457 ( .A(n298), .Y(n851) );
  INVX2TS U458 ( .A(writeIn[43]), .Y(n299) );
  INVX2TS U459 ( .A(n299), .Y(n852) );
  INVX2TS U460 ( .A(n299), .Y(n853) );
  INVX2TS U461 ( .A(writeIn[44]), .Y(n300) );
  INVX2TS U462 ( .A(n300), .Y(n854) );
  INVX2TS U463 ( .A(n300), .Y(n855) );
  INVX2TS U464 ( .A(writeIn[45]), .Y(n301) );
  INVX2TS U465 ( .A(n301), .Y(n856) );
  INVX2TS U466 ( .A(n301), .Y(n857) );
  INVX2TS U467 ( .A(writeIn[46]), .Y(n302) );
  INVX2TS U468 ( .A(n302), .Y(n858) );
  INVX2TS U469 ( .A(n302), .Y(n859) );
  INVX2TS U470 ( .A(writeIn[47]), .Y(n303) );
  INVX2TS U471 ( .A(n303), .Y(n860) );
  INVX2TS U472 ( .A(n303), .Y(n861) );
  INVX2TS U473 ( .A(writeIn[48]), .Y(n304) );
  INVX2TS U474 ( .A(n304), .Y(n862) );
  INVX2TS U475 ( .A(n304), .Y(n863) );
  INVX2TS U476 ( .A(writeIn[49]), .Y(n305) );
  INVX2TS U477 ( .A(n305), .Y(n864) );
  INVX2TS U478 ( .A(n305), .Y(n865) );
  INVX2TS U479 ( .A(writeIn[50]), .Y(n306) );
  INVX2TS U480 ( .A(n306), .Y(n866) );
  INVX2TS U481 ( .A(n306), .Y(n867) );
  INVX2TS U482 ( .A(writeIn[51]), .Y(n307) );
  INVX2TS U483 ( .A(n307), .Y(n868) );
  INVX2TS U484 ( .A(n307), .Y(n869) );
  INVX2TS U485 ( .A(writeIn[52]), .Y(n308) );
  INVX2TS U486 ( .A(n308), .Y(n870) );
  INVX2TS U487 ( .A(n308), .Y(n871) );
  INVX2TS U488 ( .A(writeIn[53]), .Y(n309) );
  INVX2TS U489 ( .A(n309), .Y(n872) );
  INVX2TS U490 ( .A(n309), .Y(n873) );
  INVX2TS U491 ( .A(writeIn[54]), .Y(n310) );
  INVX2TS U492 ( .A(n310), .Y(n874) );
  INVX2TS U493 ( .A(n310), .Y(n875) );
  INVX2TS U494 ( .A(writeIn[55]), .Y(n311) );
  INVX2TS U495 ( .A(n311), .Y(n876) );
  INVX2TS U496 ( .A(n311), .Y(n877) );
  INVX2TS U497 ( .A(writeIn[56]), .Y(n312) );
  INVX2TS U498 ( .A(n312), .Y(n878) );
  INVX2TS U499 ( .A(n312), .Y(n879) );
  INVX2TS U500 ( .A(writeIn[57]), .Y(n313) );
  INVX2TS U501 ( .A(n313), .Y(n880) );
  INVX2TS U502 ( .A(n313), .Y(n881) );
  INVX2TS U503 ( .A(writeIn[58]), .Y(n314) );
  INVX2TS U504 ( .A(n314), .Y(n882) );
  INVX2TS U505 ( .A(n314), .Y(n883) );
  INVX2TS U506 ( .A(writeIn[59]), .Y(n315) );
  INVX2TS U507 ( .A(n315), .Y(n884) );
  INVX2TS U508 ( .A(n315), .Y(n885) );
  INVX2TS U509 ( .A(NodeSelect[2]), .Y(n318) );
  INVX2TS U510 ( .A(n318), .Y(n336) );
  INVX2TS U511 ( .A(NodeSelect[0]), .Y(n323) );
  INVX2TS U512 ( .A(n323), .Y(n320) );
  INVX2TS U513 ( .A(NodeSelect[1]), .Y(n330) );
  INVX2TS U514 ( .A(n330), .Y(n333) );
  NAND2X1TS U515 ( .A(n320), .B(n333), .Y(n316) );
  NOR2XLTS U516 ( .A(n336), .B(n316), .Y(n600) );
  CLKBUFX2TS U517 ( .A(n600), .Y(n711) );
  CLKBUFX2TS U518 ( .A(n711), .Y(n402) );
  INVX2TS U519 ( .A(writeEnable), .Y(n331) );
  INVX2TS U520 ( .A(n331), .Y(n325) );
  NOR2BX1TS U521 ( .AN(n402), .B(n331), .Y(n327) );
  CLKBUFX2TS U522 ( .A(n327), .Y(n354) );
  CLKBUFX2TS U523 ( .A(n354), .Y(n317) );
  CLKBUFX2TS U524 ( .A(n317), .Y(n951) );
  CLKBUFX2TS U525 ( .A(n317), .Y(n950) );
  CLKBUFX2TS U526 ( .A(n317), .Y(n949) );
  CLKBUFX2TS U527 ( .A(n317), .Y(n947) );
  INVX2TS U528 ( .A(n318), .Y(n339) );
  NOR3XLTS U529 ( .A(n320), .B(n332), .C(n324), .Y(n599) );
  CLKBUFX2TS U530 ( .A(n599), .Y(n709) );
  CLKBUFX2TS U531 ( .A(n709), .Y(n400) );
  CLKAND2X2TS U532 ( .A(n400), .B(n325), .Y(n348) );
  CLKBUFX2TS U533 ( .A(n348), .Y(n898) );
  CLKBUFX2TS U534 ( .A(n348), .Y(n326) );
  CLKBUFX2TS U535 ( .A(n326), .Y(n319) );
  CLKBUFX2TS U536 ( .A(n319), .Y(n993) );
  CLKBUFX2TS U537 ( .A(n319), .Y(n992) );
  CLKBUFX2TS U538 ( .A(n319), .Y(n991) );
  CLKBUFX2TS U539 ( .A(n319), .Y(n990) );
  NOR3XLTS U540 ( .A(n332), .B(n337), .C(n324), .Y(n601) );
  CLKBUFX2TS U541 ( .A(n601), .Y(n713) );
  CLKBUFX2TS U542 ( .A(n713), .Y(n404) );
  NOR2BX1TS U543 ( .AN(n404), .B(n331), .Y(n321) );
  CLKBUFX2TS U544 ( .A(n321), .Y(n900) );
  CLKBUFX2TS U545 ( .A(n321), .Y(n358) );
  CLKBUFX2TS U546 ( .A(n358), .Y(n322) );
  CLKBUFX2TS U547 ( .A(n322), .Y(n1006) );
  CLKBUFX2TS U548 ( .A(n322), .Y(n1005) );
  CLKBUFX2TS U549 ( .A(n322), .Y(n1004) );
  CLKBUFX2TS U550 ( .A(n322), .Y(n1002) );
  INVX2TS U551 ( .A(n323), .Y(n335) );
  NOR3XLTS U552 ( .A(n336), .B(n335), .C(n324), .Y(n598) );
  CLKBUFX2TS U553 ( .A(n598), .Y(n707) );
  CLKBUFX2TS U554 ( .A(n707), .Y(n398) );
  CLKAND2X2TS U555 ( .A(n398), .B(n325), .Y(n349) );
  CLKBUFX2TS U556 ( .A(n349), .Y(n328) );
  CLKBUFX2TS U557 ( .A(n328), .Y(n933) );
  CLKBUFX2TS U558 ( .A(n328), .Y(n931) );
  CLKBUFX2TS U559 ( .A(n328), .Y(n930) );
  CLKBUFX2TS U560 ( .A(n354), .Y(n948) );
  CLKBUFX2TS U561 ( .A(n326), .Y(n988) );
  CLKBUFX2TS U562 ( .A(n326), .Y(n986) );
  CLKBUFX2TS U563 ( .A(n326), .Y(n985) );
  CLKBUFX2TS U564 ( .A(n358), .Y(n1003) );
  CLKBUFX2TS U565 ( .A(n349), .Y(n890) );
  CLKBUFX2TS U566 ( .A(n890), .Y(n891) );
  CLKBUFX2TS U567 ( .A(n891), .Y(n943) );
  CLKBUFX2TS U568 ( .A(n891), .Y(n942) );
  CLKBUFX2TS U569 ( .A(n327), .Y(n892) );
  CLKBUFX2TS U570 ( .A(n892), .Y(n893) );
  CLKBUFX2TS U571 ( .A(n893), .Y(n956) );
  CLKBUFX2TS U572 ( .A(n893), .Y(n955) );
  CLKBUFX2TS U573 ( .A(n898), .Y(n899) );
  CLKBUFX2TS U574 ( .A(n899), .Y(n997) );
  CLKBUFX2TS U575 ( .A(n900), .Y(n901) );
  CLKBUFX2TS U576 ( .A(n901), .Y(n1011) );
  CLKBUFX2TS U577 ( .A(n901), .Y(n1010) );
  CLKBUFX2TS U578 ( .A(n328), .Y(n329) );
  CLKBUFX2TS U579 ( .A(n329), .Y(n938) );
  CLKBUFX2TS U580 ( .A(n329), .Y(n937) );
  CLKBUFX2TS U581 ( .A(n329), .Y(n936) );
  CLKBUFX2TS U582 ( .A(n329), .Y(n935) );
  CLKBUFX2TS U583 ( .A(n899), .Y(n998) );
  INVX2TS U584 ( .A(n330), .Y(n338) );
  NOR3XLTS U585 ( .A(n335), .B(n338), .C(n332), .Y(n415) );
  CLKBUFX2TS U586 ( .A(n415), .Y(n443) );
  CLKBUFX2TS U587 ( .A(n443), .Y(n401) );
  INVX2TS U588 ( .A(n331), .Y(n340) );
  CLKAND2X2TS U589 ( .A(n401), .B(n340), .Y(n352) );
  CLKBUFX2TS U590 ( .A(n352), .Y(n341) );
  CLKBUFX2TS U591 ( .A(n341), .Y(n342) );
  CLKBUFX2TS U592 ( .A(n342), .Y(n963) );
  CLKBUFX2TS U593 ( .A(n342), .Y(n962) );
  NOR3XLTS U594 ( .A(n333), .B(n337), .C(n332), .Y(n417) );
  CLKBUFX2TS U595 ( .A(n417), .Y(n445) );
  CLKBUFX2TS U596 ( .A(n445), .Y(n405) );
  CLKAND2X2TS U597 ( .A(n405), .B(n340), .Y(n353) );
  CLKBUFX2TS U598 ( .A(n353), .Y(n347) );
  CLKBUFX2TS U599 ( .A(n347), .Y(n334) );
  CLKBUFX2TS U600 ( .A(n334), .Y(n979) );
  CLKBUFX2TS U601 ( .A(n334), .Y(n978) );
  CLKBUFX2TS U602 ( .A(n334), .Y(n977) );
  CLKBUFX2TS U603 ( .A(n334), .Y(n976) );
  NOR3XLTS U604 ( .A(n336), .B(n335), .C(n338), .Y(n414) );
  CLKBUFX2TS U605 ( .A(n414), .Y(n442) );
  CLKBUFX2TS U606 ( .A(n442), .Y(n399) );
  CLKAND2X2TS U607 ( .A(n399), .B(n340), .Y(n350) );
  CLKBUFX2TS U608 ( .A(n350), .Y(n886) );
  CLKBUFX2TS U609 ( .A(n886), .Y(n887) );
  CLKBUFX2TS U610 ( .A(n887), .Y(n915) );
  CLKBUFX2TS U611 ( .A(n887), .Y(n914) );
  NOR3XLTS U612 ( .A(n339), .B(n338), .C(n337), .Y(n416) );
  CLKBUFX2TS U613 ( .A(n416), .Y(n444) );
  CLKBUFX2TS U614 ( .A(n444), .Y(n403) );
  CLKAND2X2TS U615 ( .A(n403), .B(n340), .Y(n351) );
  CLKBUFX2TS U616 ( .A(n351), .Y(n888) );
  CLKBUFX2TS U617 ( .A(n888), .Y(n889) );
  CLKBUFX2TS U618 ( .A(n889), .Y(n929) );
  CLKBUFX2TS U619 ( .A(n889), .Y(n928) );
  CLKBUFX2TS U620 ( .A(n352), .Y(n894) );
  CLKBUFX2TS U621 ( .A(n894), .Y(n895) );
  CLKBUFX2TS U622 ( .A(n895), .Y(n970) );
  CLKBUFX2TS U623 ( .A(n895), .Y(n969) );
  CLKBUFX2TS U624 ( .A(n353), .Y(n896) );
  CLKBUFX2TS U625 ( .A(n896), .Y(n897) );
  CLKBUFX2TS U626 ( .A(n897), .Y(n984) );
  CLKBUFX2TS U627 ( .A(n897), .Y(n983) );
  CLKBUFX2TS U628 ( .A(n350), .Y(n345) );
  CLKBUFX2TS U629 ( .A(n345), .Y(n905) );
  CLKBUFX2TS U630 ( .A(n345), .Y(n903) );
  CLKBUFX2TS U631 ( .A(n345), .Y(n902) );
  CLKBUFX2TS U632 ( .A(n351), .Y(n343) );
  CLKBUFX2TS U633 ( .A(n343), .Y(n919) );
  CLKBUFX2TS U634 ( .A(n343), .Y(n917) );
  CLKBUFX2TS U635 ( .A(n343), .Y(n916) );
  CLKBUFX2TS U636 ( .A(n341), .Y(n960) );
  CLKBUFX2TS U637 ( .A(n341), .Y(n958) );
  CLKBUFX2TS U638 ( .A(n341), .Y(n957) );
  CLKBUFX2TS U639 ( .A(n342), .Y(n964) );
  CLKBUFX2TS U640 ( .A(n342), .Y(n965) );
  CLKBUFX2TS U641 ( .A(n343), .Y(n344) );
  CLKBUFX2TS U642 ( .A(n344), .Y(n921) );
  CLKBUFX2TS U643 ( .A(n344), .Y(n922) );
  CLKBUFX2TS U644 ( .A(n344), .Y(n923) );
  CLKBUFX2TS U645 ( .A(n344), .Y(n924) );
  CLKBUFX2TS U646 ( .A(n345), .Y(n346) );
  CLKBUFX2TS U647 ( .A(n346), .Y(n907) );
  CLKBUFX2TS U648 ( .A(n346), .Y(n908) );
  CLKBUFX2TS U649 ( .A(n346), .Y(n909) );
  CLKBUFX2TS U650 ( .A(n346), .Y(n910) );
  CLKBUFX2TS U651 ( .A(n347), .Y(n971) );
  CLKBUFX2TS U652 ( .A(n347), .Y(n972) );
  CLKBUFX2TS U653 ( .A(n347), .Y(n974) );
  CLKBUFX2TS U654 ( .A(n349), .Y(n932) );
  CLKBUFX2TS U655 ( .A(n348), .Y(n989) );
  CLKBUFX2TS U656 ( .A(n348), .Y(n987) );
  CLKBUFX2TS U657 ( .A(n349), .Y(n934) );
  CLKBUFX2TS U658 ( .A(n350), .Y(n906) );
  CLKBUFX2TS U659 ( .A(n350), .Y(n904) );
  CLKBUFX2TS U660 ( .A(n351), .Y(n920) );
  CLKBUFX2TS U661 ( .A(n351), .Y(n918) );
  CLKBUFX2TS U662 ( .A(n352), .Y(n961) );
  CLKBUFX2TS U663 ( .A(n352), .Y(n959) );
  CLKBUFX2TS U664 ( .A(n353), .Y(n973) );
  CLKBUFX2TS U665 ( .A(n353), .Y(n975) );
  CLKBUFX2TS U666 ( .A(n892), .Y(n361) );
  CLKBUFX2TS U667 ( .A(n361), .Y(n952) );
  CLKBUFX2TS U668 ( .A(n354), .Y(n355) );
  CLKBUFX2TS U669 ( .A(n355), .Y(n946) );
  CLKBUFX2TS U670 ( .A(n355), .Y(n945) );
  CLKBUFX2TS U671 ( .A(n355), .Y(n944) );
  CLKBUFX2TS U672 ( .A(n898), .Y(n356) );
  CLKBUFX2TS U673 ( .A(n356), .Y(n996) );
  CLKBUFX2TS U674 ( .A(n356), .Y(n995) );
  CLKBUFX2TS U675 ( .A(n356), .Y(n994) );
  CLKBUFX2TS U676 ( .A(n361), .Y(n953) );
  CLKBUFX2TS U677 ( .A(n900), .Y(n357) );
  CLKBUFX2TS U678 ( .A(n357), .Y(n1009) );
  CLKBUFX2TS U679 ( .A(n357), .Y(n1008) );
  CLKBUFX2TS U680 ( .A(n357), .Y(n1007) );
  CLKBUFX2TS U681 ( .A(n358), .Y(n359) );
  CLKBUFX2TS U682 ( .A(n359), .Y(n1001) );
  CLKBUFX2TS U683 ( .A(n359), .Y(n1000) );
  CLKBUFX2TS U684 ( .A(n359), .Y(n999) );
  CLKBUFX2TS U685 ( .A(n890), .Y(n360) );
  CLKBUFX2TS U686 ( .A(n360), .Y(n941) );
  CLKBUFX2TS U687 ( .A(n360), .Y(n940) );
  CLKBUFX2TS U688 ( .A(n360), .Y(n939) );
  CLKBUFX2TS U689 ( .A(n361), .Y(n954) );
  CLKBUFX2TS U690 ( .A(n886), .Y(n362) );
  CLKBUFX2TS U691 ( .A(n362), .Y(n913) );
  CLKBUFX2TS U692 ( .A(n362), .Y(n912) );
  CLKBUFX2TS U693 ( .A(n362), .Y(n911) );
  CLKBUFX2TS U694 ( .A(n888), .Y(n363) );
  CLKBUFX2TS U695 ( .A(n363), .Y(n927) );
  CLKBUFX2TS U696 ( .A(n363), .Y(n926) );
  CLKBUFX2TS U697 ( .A(n363), .Y(n925) );
  CLKBUFX2TS U698 ( .A(n894), .Y(n364) );
  CLKBUFX2TS U699 ( .A(n364), .Y(n968) );
  CLKBUFX2TS U700 ( .A(n364), .Y(n967) );
  CLKBUFX2TS U701 ( .A(n364), .Y(n966) );
  CLKBUFX2TS U702 ( .A(n896), .Y(n365) );
  CLKBUFX2TS U703 ( .A(n365), .Y(n982) );
  CLKBUFX2TS U704 ( .A(n365), .Y(n981) );
  CLKBUFX2TS U705 ( .A(n365), .Y(n980) );
  CLKBUFX2TS U706 ( .A(n442), .Y(n379) );
  CLKBUFX2TS U707 ( .A(n707), .Y(n378) );
  AOI22X1TS U708 ( .A0(n379), .A1(readOutBus[59]), .B0(n378), .B1(
        readOutBus[179]), .Y(n369) );
  CLKBUFX2TS U709 ( .A(n443), .Y(n381) );
  CLKBUFX2TS U710 ( .A(n709), .Y(n380) );
  AOI22X1TS U711 ( .A0(n381), .A1(readOutBus[299]), .B0(n380), .B1(
        readOutBus[419]), .Y(n368) );
  CLKBUFX2TS U712 ( .A(n444), .Y(n383) );
  CLKBUFX2TS U713 ( .A(n711), .Y(n382) );
  AOI22X1TS U714 ( .A0(n383), .A1(readOutBus[119]), .B0(n382), .B1(
        readOutBus[239]), .Y(n367) );
  CLKBUFX2TS U715 ( .A(n445), .Y(n385) );
  CLKBUFX2TS U716 ( .A(n713), .Y(n384) );
  AOI22X1TS U717 ( .A0(n385), .A1(readOutBus[359]), .B0(n384), .B1(
        readOutBus[479]), .Y(n366) );
  NAND4XLTS U718 ( .A(n369), .B(n368), .C(n367), .D(n366), .Y(readOut[59]) );
  AOI22X1TS U719 ( .A0(n379), .A1(readOutBus[58]), .B0(n378), .B1(
        readOutBus[178]), .Y(n373) );
  AOI22X1TS U720 ( .A0(n381), .A1(readOutBus[298]), .B0(n380), .B1(
        readOutBus[418]), .Y(n372) );
  AOI22X1TS U721 ( .A0(n383), .A1(readOutBus[118]), .B0(n382), .B1(
        readOutBus[238]), .Y(n371) );
  AOI22X1TS U722 ( .A0(n385), .A1(readOutBus[358]), .B0(n384), .B1(
        readOutBus[478]), .Y(n370) );
  NAND4XLTS U723 ( .A(n373), .B(n372), .C(n371), .D(n370), .Y(readOut[58]) );
  AOI22X1TS U724 ( .A0(n379), .A1(readOutBus[57]), .B0(n378), .B1(
        readOutBus[177]), .Y(n377) );
  AOI22X1TS U725 ( .A0(n381), .A1(readOutBus[297]), .B0(n380), .B1(
        readOutBus[417]), .Y(n376) );
  AOI22X1TS U726 ( .A0(n383), .A1(readOutBus[117]), .B0(n382), .B1(
        readOutBus[237]), .Y(n375) );
  AOI22X1TS U727 ( .A0(n385), .A1(readOutBus[357]), .B0(n384), .B1(
        readOutBus[477]), .Y(n374) );
  NAND4XLTS U728 ( .A(n377), .B(n376), .C(n375), .D(n374), .Y(readOut[57]) );
  AOI22X1TS U729 ( .A0(n379), .A1(readOutBus[56]), .B0(n378), .B1(
        readOutBus[176]), .Y(n389) );
  AOI22X1TS U730 ( .A0(n381), .A1(readOutBus[296]), .B0(n380), .B1(
        readOutBus[416]), .Y(n388) );
  AOI22X1TS U731 ( .A0(n383), .A1(readOutBus[116]), .B0(n382), .B1(
        readOutBus[236]), .Y(n387) );
  AOI22X1TS U732 ( .A0(n385), .A1(readOutBus[356]), .B0(n384), .B1(
        readOutBus[476]), .Y(n386) );
  NAND4XLTS U733 ( .A(n389), .B(n388), .C(n387), .D(n386), .Y(readOut[56]) );
  AOI22X1TS U734 ( .A0(n399), .A1(readOutBus[55]), .B0(n398), .B1(
        readOutBus[175]), .Y(n393) );
  AOI22X1TS U735 ( .A0(n401), .A1(readOutBus[295]), .B0(n400), .B1(
        readOutBus[415]), .Y(n392) );
  AOI22X1TS U736 ( .A0(n403), .A1(readOutBus[115]), .B0(n402), .B1(
        readOutBus[235]), .Y(n391) );
  AOI22X1TS U737 ( .A0(n405), .A1(readOutBus[355]), .B0(n404), .B1(
        readOutBus[475]), .Y(n390) );
  NAND4XLTS U738 ( .A(n393), .B(n392), .C(n391), .D(n390), .Y(readOut[55]) );
  AOI22X1TS U739 ( .A0(n399), .A1(readOutBus[54]), .B0(n398), .B1(
        readOutBus[174]), .Y(n397) );
  AOI22X1TS U740 ( .A0(n401), .A1(readOutBus[294]), .B0(n400), .B1(
        readOutBus[414]), .Y(n396) );
  AOI22X1TS U741 ( .A0(n403), .A1(readOutBus[114]), .B0(n402), .B1(
        readOutBus[234]), .Y(n395) );
  AOI22X1TS U742 ( .A0(n405), .A1(readOutBus[354]), .B0(n404), .B1(
        readOutBus[474]), .Y(n394) );
  NAND4XLTS U743 ( .A(n397), .B(n396), .C(n395), .D(n394), .Y(readOut[54]) );
  AOI22X1TS U744 ( .A0(n399), .A1(readOutBus[53]), .B0(n398), .B1(
        readOutBus[173]), .Y(n409) );
  AOI22X1TS U745 ( .A0(n401), .A1(readOutBus[293]), .B0(n400), .B1(
        readOutBus[413]), .Y(n408) );
  AOI22X1TS U746 ( .A0(n403), .A1(readOutBus[113]), .B0(n402), .B1(
        readOutBus[233]), .Y(n407) );
  AOI22X1TS U747 ( .A0(n405), .A1(readOutBus[353]), .B0(n404), .B1(
        readOutBus[473]), .Y(n406) );
  NAND4XLTS U748 ( .A(n409), .B(n408), .C(n407), .D(n406), .Y(readOut[53]) );
  AOI22X1TS U749 ( .A0(n442), .A1(readOutBus[52]), .B0(n707), .B1(
        readOutBus[172]), .Y(n413) );
  AOI22X1TS U750 ( .A0(n443), .A1(readOutBus[292]), .B0(n709), .B1(
        readOutBus[412]), .Y(n412) );
  AOI22X1TS U751 ( .A0(n444), .A1(readOutBus[112]), .B0(n711), .B1(
        readOutBus[232]), .Y(n411) );
  AOI22X1TS U752 ( .A0(n445), .A1(readOutBus[352]), .B0(n713), .B1(
        readOutBus[472]), .Y(n410) );
  NAND4XLTS U753 ( .A(n413), .B(n412), .C(n411), .D(n410), .Y(readOut[52]) );
  CLKBUFX2TS U754 ( .A(n414), .Y(n626) );
  CLKBUFX2TS U755 ( .A(n626), .Y(n431) );
  CLKBUFX2TS U756 ( .A(n598), .Y(n627) );
  CLKBUFX2TS U757 ( .A(n627), .Y(n578) );
  CLKBUFX2TS U758 ( .A(n578), .Y(n430) );
  AOI22X1TS U759 ( .A0(n431), .A1(readOutBus[51]), .B0(n430), .B1(
        readOutBus[171]), .Y(n421) );
  CLKBUFX2TS U760 ( .A(n415), .Y(n628) );
  CLKBUFX2TS U761 ( .A(n628), .Y(n433) );
  CLKBUFX2TS U762 ( .A(n599), .Y(n629) );
  CLKBUFX2TS U763 ( .A(n629), .Y(n579) );
  CLKBUFX2TS U764 ( .A(n579), .Y(n432) );
  AOI22X1TS U765 ( .A0(n433), .A1(readOutBus[291]), .B0(n432), .B1(
        readOutBus[411]), .Y(n420) );
  CLKBUFX2TS U766 ( .A(n416), .Y(n630) );
  CLKBUFX2TS U767 ( .A(n630), .Y(n435) );
  CLKBUFX2TS U768 ( .A(n600), .Y(n580) );
  CLKBUFX2TS U769 ( .A(n580), .Y(n434) );
  AOI22X1TS U770 ( .A0(n435), .A1(readOutBus[111]), .B0(n434), .B1(
        readOutBus[231]), .Y(n419) );
  CLKBUFX2TS U771 ( .A(n417), .Y(n632) );
  CLKBUFX2TS U772 ( .A(n632), .Y(n437) );
  CLKBUFX2TS U773 ( .A(n601), .Y(n633) );
  CLKBUFX2TS U774 ( .A(n633), .Y(n581) );
  CLKBUFX2TS U775 ( .A(n581), .Y(n436) );
  AOI22X1TS U776 ( .A0(n437), .A1(readOutBus[351]), .B0(n436), .B1(
        readOutBus[471]), .Y(n418) );
  NAND4XLTS U777 ( .A(n421), .B(n420), .C(n419), .D(n418), .Y(readOut[51]) );
  AOI22X1TS U778 ( .A0(n431), .A1(readOutBus[50]), .B0(n430), .B1(
        readOutBus[170]), .Y(n425) );
  AOI22X1TS U779 ( .A0(n433), .A1(readOutBus[290]), .B0(n432), .B1(
        readOutBus[410]), .Y(n424) );
  AOI22X1TS U780 ( .A0(n435), .A1(readOutBus[110]), .B0(n434), .B1(
        readOutBus[230]), .Y(n423) );
  AOI22X1TS U781 ( .A0(n437), .A1(readOutBus[350]), .B0(n436), .B1(
        readOutBus[470]), .Y(n422) );
  NAND4XLTS U782 ( .A(n425), .B(n424), .C(n423), .D(n422), .Y(readOut[50]) );
  AOI22X1TS U783 ( .A0(n431), .A1(readOutBus[49]), .B0(n430), .B1(
        readOutBus[169]), .Y(n429) );
  AOI22X1TS U784 ( .A0(n433), .A1(readOutBus[289]), .B0(n432), .B1(
        readOutBus[409]), .Y(n428) );
  AOI22X1TS U785 ( .A0(n435), .A1(readOutBus[109]), .B0(n434), .B1(
        readOutBus[229]), .Y(n427) );
  AOI22X1TS U786 ( .A0(n437), .A1(readOutBus[349]), .B0(n436), .B1(
        readOutBus[469]), .Y(n426) );
  NAND4XLTS U787 ( .A(n429), .B(n428), .C(n427), .D(n426), .Y(readOut[49]) );
  AOI22X1TS U788 ( .A0(n431), .A1(readOutBus[48]), .B0(n430), .B1(
        readOutBus[168]), .Y(n441) );
  AOI22X1TS U789 ( .A0(n433), .A1(readOutBus[288]), .B0(n432), .B1(
        readOutBus[408]), .Y(n440) );
  AOI22X1TS U790 ( .A0(n435), .A1(readOutBus[108]), .B0(n434), .B1(
        readOutBus[228]), .Y(n439) );
  AOI22X1TS U791 ( .A0(n437), .A1(readOutBus[348]), .B0(n436), .B1(
        readOutBus[468]), .Y(n438) );
  NAND4XLTS U792 ( .A(n441), .B(n440), .C(n439), .D(n438), .Y(readOut[48]) );
  CLKBUFX2TS U793 ( .A(n442), .Y(n459) );
  CLKBUFX2TS U794 ( .A(n578), .Y(n458) );
  AOI22X1TS U795 ( .A0(n459), .A1(readOutBus[47]), .B0(n458), .B1(
        readOutBus[167]), .Y(n449) );
  CLKBUFX2TS U796 ( .A(n443), .Y(n461) );
  CLKBUFX2TS U797 ( .A(n579), .Y(n460) );
  AOI22X1TS U798 ( .A0(n461), .A1(readOutBus[287]), .B0(n460), .B1(
        readOutBus[407]), .Y(n448) );
  CLKBUFX2TS U799 ( .A(n444), .Y(n463) );
  CLKBUFX2TS U800 ( .A(n580), .Y(n462) );
  AOI22X1TS U801 ( .A0(n463), .A1(readOutBus[107]), .B0(n462), .B1(
        readOutBus[227]), .Y(n447) );
  CLKBUFX2TS U802 ( .A(n445), .Y(n465) );
  CLKBUFX2TS U803 ( .A(n581), .Y(n464) );
  AOI22X1TS U804 ( .A0(n465), .A1(readOutBus[347]), .B0(n464), .B1(
        readOutBus[467]), .Y(n446) );
  NAND4XLTS U805 ( .A(n449), .B(n448), .C(n447), .D(n446), .Y(readOut[47]) );
  AOI22X1TS U806 ( .A0(n459), .A1(readOutBus[46]), .B0(n458), .B1(
        readOutBus[166]), .Y(n453) );
  AOI22X1TS U807 ( .A0(n461), .A1(readOutBus[286]), .B0(n460), .B1(
        readOutBus[406]), .Y(n452) );
  AOI22X1TS U808 ( .A0(n463), .A1(readOutBus[106]), .B0(n462), .B1(
        readOutBus[226]), .Y(n451) );
  AOI22X1TS U809 ( .A0(n465), .A1(readOutBus[346]), .B0(n464), .B1(
        readOutBus[466]), .Y(n450) );
  NAND4XLTS U810 ( .A(n453), .B(n452), .C(n451), .D(n450), .Y(readOut[46]) );
  AOI22X1TS U811 ( .A0(n459), .A1(readOutBus[45]), .B0(n458), .B1(
        readOutBus[165]), .Y(n457) );
  AOI22X1TS U812 ( .A0(n461), .A1(readOutBus[285]), .B0(n460), .B1(
        readOutBus[405]), .Y(n456) );
  AOI22X1TS U813 ( .A0(n463), .A1(readOutBus[105]), .B0(n462), .B1(
        readOutBus[225]), .Y(n455) );
  AOI22X1TS U814 ( .A0(n465), .A1(readOutBus[345]), .B0(n464), .B1(
        readOutBus[465]), .Y(n454) );
  NAND4XLTS U815 ( .A(n457), .B(n456), .C(n455), .D(n454), .Y(readOut[45]) );
  AOI22X1TS U816 ( .A0(n459), .A1(readOutBus[44]), .B0(n458), .B1(
        readOutBus[164]), .Y(n469) );
  AOI22X1TS U817 ( .A0(n461), .A1(readOutBus[284]), .B0(n460), .B1(
        readOutBus[404]), .Y(n468) );
  AOI22X1TS U818 ( .A0(n463), .A1(readOutBus[104]), .B0(n462), .B1(
        readOutBus[224]), .Y(n467) );
  AOI22X1TS U819 ( .A0(n465), .A1(readOutBus[344]), .B0(n464), .B1(
        readOutBus[464]), .Y(n466) );
  NAND4XLTS U820 ( .A(n469), .B(n468), .C(n467), .D(n466), .Y(readOut[44]) );
  CLKBUFX2TS U821 ( .A(n626), .Y(n734) );
  CLKBUFX2TS U822 ( .A(n734), .Y(n483) );
  CLKBUFX2TS U823 ( .A(n578), .Y(n482) );
  AOI22X1TS U824 ( .A0(n483), .A1(readOutBus[43]), .B0(n482), .B1(
        readOutBus[163]), .Y(n473) );
  CLKBUFX2TS U825 ( .A(n628), .Y(n736) );
  CLKBUFX2TS U826 ( .A(n736), .Y(n485) );
  CLKBUFX2TS U827 ( .A(n579), .Y(n484) );
  AOI22X1TS U828 ( .A0(n485), .A1(readOutBus[283]), .B0(n484), .B1(
        readOutBus[403]), .Y(n472) );
  CLKBUFX2TS U829 ( .A(n630), .Y(n738) );
  CLKBUFX2TS U830 ( .A(n738), .Y(n487) );
  CLKBUFX2TS U831 ( .A(n580), .Y(n486) );
  AOI22X1TS U832 ( .A0(n487), .A1(readOutBus[103]), .B0(n486), .B1(
        readOutBus[223]), .Y(n471) );
  CLKBUFX2TS U833 ( .A(n632), .Y(n740) );
  CLKBUFX2TS U834 ( .A(n740), .Y(n489) );
  CLKBUFX2TS U835 ( .A(n581), .Y(n488) );
  AOI22X1TS U836 ( .A0(n489), .A1(readOutBus[343]), .B0(n488), .B1(
        readOutBus[463]), .Y(n470) );
  NAND4XLTS U837 ( .A(n473), .B(n472), .C(n471), .D(n470), .Y(readOut[43]) );
  AOI22X1TS U838 ( .A0(n483), .A1(readOutBus[42]), .B0(n482), .B1(
        readOutBus[162]), .Y(n477) );
  AOI22X1TS U839 ( .A0(n485), .A1(readOutBus[282]), .B0(n484), .B1(
        readOutBus[402]), .Y(n476) );
  AOI22X1TS U840 ( .A0(n487), .A1(readOutBus[102]), .B0(n486), .B1(
        readOutBus[222]), .Y(n475) );
  AOI22X1TS U841 ( .A0(n489), .A1(readOutBus[342]), .B0(n488), .B1(
        readOutBus[462]), .Y(n474) );
  NAND4XLTS U842 ( .A(n477), .B(n476), .C(n475), .D(n474), .Y(readOut[42]) );
  AOI22X1TS U843 ( .A0(n483), .A1(readOutBus[41]), .B0(n482), .B1(
        readOutBus[161]), .Y(n481) );
  AOI22X1TS U844 ( .A0(n485), .A1(readOutBus[281]), .B0(n484), .B1(
        readOutBus[401]), .Y(n480) );
  AOI22X1TS U845 ( .A0(n487), .A1(readOutBus[101]), .B0(n486), .B1(
        readOutBus[221]), .Y(n479) );
  AOI22X1TS U846 ( .A0(n489), .A1(readOutBus[341]), .B0(n488), .B1(
        readOutBus[461]), .Y(n478) );
  NAND4XLTS U847 ( .A(n481), .B(n480), .C(n479), .D(n478), .Y(readOut[41]) );
  AOI22X1TS U848 ( .A0(n483), .A1(readOutBus[40]), .B0(n482), .B1(
        readOutBus[160]), .Y(n493) );
  AOI22X1TS U849 ( .A0(n485), .A1(readOutBus[280]), .B0(n484), .B1(
        readOutBus[400]), .Y(n492) );
  AOI22X1TS U850 ( .A0(n487), .A1(readOutBus[100]), .B0(n486), .B1(
        readOutBus[220]), .Y(n491) );
  AOI22X1TS U851 ( .A0(n489), .A1(readOutBus[340]), .B0(n488), .B1(
        readOutBus[460]), .Y(n490) );
  NAND4XLTS U852 ( .A(n493), .B(n492), .C(n491), .D(n490), .Y(readOut[40]) );
  CLKBUFX2TS U853 ( .A(n734), .Y(n706) );
  CLKBUFX2TS U854 ( .A(n706), .Y(n542) );
  CLKBUFX2TS U855 ( .A(n542), .Y(n507) );
  CLKBUFX2TS U856 ( .A(n627), .Y(n586) );
  CLKBUFX2TS U857 ( .A(n586), .Y(n506) );
  AOI22X1TS U858 ( .A0(n507), .A1(readOutBus[39]), .B0(n506), .B1(
        readOutBus[159]), .Y(n497) );
  CLKBUFX2TS U859 ( .A(n736), .Y(n708) );
  CLKBUFX2TS U860 ( .A(n708), .Y(n543) );
  CLKBUFX2TS U861 ( .A(n543), .Y(n509) );
  CLKBUFX2TS U862 ( .A(n629), .Y(n588) );
  CLKBUFX2TS U863 ( .A(n588), .Y(n508) );
  AOI22X1TS U864 ( .A0(n509), .A1(readOutBus[279]), .B0(n508), .B1(
        readOutBus[399]), .Y(n496) );
  CLKBUFX2TS U865 ( .A(n738), .Y(n710) );
  CLKBUFX2TS U866 ( .A(n710), .Y(n544) );
  CLKBUFX2TS U867 ( .A(n544), .Y(n511) );
  CLKBUFX2TS U868 ( .A(n600), .Y(n631) );
  CLKBUFX2TS U869 ( .A(n631), .Y(n590) );
  CLKBUFX2TS U870 ( .A(n590), .Y(n510) );
  AOI22X1TS U871 ( .A0(n511), .A1(readOutBus[99]), .B0(n510), .B1(
        readOutBus[219]), .Y(n495) );
  CLKBUFX2TS U872 ( .A(n740), .Y(n712) );
  CLKBUFX2TS U873 ( .A(n712), .Y(n545) );
  CLKBUFX2TS U874 ( .A(n545), .Y(n513) );
  CLKBUFX2TS U875 ( .A(n633), .Y(n592) );
  CLKBUFX2TS U876 ( .A(n592), .Y(n512) );
  AOI22X1TS U877 ( .A0(n513), .A1(readOutBus[339]), .B0(n512), .B1(
        readOutBus[459]), .Y(n494) );
  NAND4XLTS U878 ( .A(n497), .B(n496), .C(n495), .D(n494), .Y(readOut[39]) );
  AOI22X1TS U879 ( .A0(n507), .A1(readOutBus[38]), .B0(n506), .B1(
        readOutBus[158]), .Y(n501) );
  AOI22X1TS U880 ( .A0(n509), .A1(readOutBus[278]), .B0(n508), .B1(
        readOutBus[398]), .Y(n500) );
  AOI22X1TS U881 ( .A0(n511), .A1(readOutBus[98]), .B0(n510), .B1(
        readOutBus[218]), .Y(n499) );
  AOI22X1TS U882 ( .A0(n513), .A1(readOutBus[338]), .B0(n512), .B1(
        readOutBus[458]), .Y(n498) );
  NAND4XLTS U883 ( .A(n501), .B(n500), .C(n499), .D(n498), .Y(readOut[38]) );
  AOI22X1TS U884 ( .A0(n507), .A1(readOutBus[37]), .B0(n506), .B1(
        readOutBus[157]), .Y(n505) );
  AOI22X1TS U885 ( .A0(n509), .A1(readOutBus[277]), .B0(n508), .B1(
        readOutBus[397]), .Y(n504) );
  AOI22X1TS U886 ( .A0(n511), .A1(readOutBus[97]), .B0(n510), .B1(
        readOutBus[217]), .Y(n503) );
  AOI22X1TS U887 ( .A0(n513), .A1(readOutBus[337]), .B0(n512), .B1(
        readOutBus[457]), .Y(n502) );
  NAND4XLTS U888 ( .A(n505), .B(n504), .C(n503), .D(n502), .Y(readOut[37]) );
  AOI22X1TS U889 ( .A0(n507), .A1(readOutBus[36]), .B0(n506), .B1(
        readOutBus[156]), .Y(n517) );
  AOI22X1TS U890 ( .A0(n509), .A1(readOutBus[276]), .B0(n508), .B1(
        readOutBus[396]), .Y(n516) );
  AOI22X1TS U891 ( .A0(n511), .A1(readOutBus[96]), .B0(n510), .B1(
        readOutBus[216]), .Y(n515) );
  AOI22X1TS U892 ( .A0(n513), .A1(readOutBus[336]), .B0(n512), .B1(
        readOutBus[456]), .Y(n514) );
  NAND4XLTS U893 ( .A(n517), .B(n516), .C(n515), .D(n514), .Y(readOut[36]) );
  CLKBUFX2TS U894 ( .A(n542), .Y(n531) );
  CLKBUFX2TS U895 ( .A(n586), .Y(n530) );
  AOI22X1TS U896 ( .A0(n531), .A1(readOutBus[35]), .B0(n530), .B1(
        readOutBus[155]), .Y(n521) );
  CLKBUFX2TS U897 ( .A(n543), .Y(n533) );
  CLKBUFX2TS U898 ( .A(n588), .Y(n532) );
  AOI22X1TS U899 ( .A0(n533), .A1(readOutBus[275]), .B0(n532), .B1(
        readOutBus[395]), .Y(n520) );
  CLKBUFX2TS U900 ( .A(n544), .Y(n535) );
  CLKBUFX2TS U901 ( .A(n590), .Y(n534) );
  AOI22X1TS U902 ( .A0(n535), .A1(readOutBus[95]), .B0(n534), .B1(
        readOutBus[215]), .Y(n519) );
  CLKBUFX2TS U903 ( .A(n545), .Y(n537) );
  CLKBUFX2TS U904 ( .A(n592), .Y(n536) );
  AOI22X1TS U905 ( .A0(n537), .A1(readOutBus[335]), .B0(n536), .B1(
        readOutBus[455]), .Y(n518) );
  NAND4XLTS U906 ( .A(n521), .B(n520), .C(n519), .D(n518), .Y(readOut[35]) );
  AOI22X1TS U907 ( .A0(n531), .A1(readOutBus[34]), .B0(n530), .B1(
        readOutBus[154]), .Y(n525) );
  AOI22X1TS U908 ( .A0(n533), .A1(readOutBus[274]), .B0(n532), .B1(
        readOutBus[394]), .Y(n524) );
  AOI22X1TS U909 ( .A0(n535), .A1(readOutBus[94]), .B0(n534), .B1(
        readOutBus[214]), .Y(n523) );
  AOI22X1TS U910 ( .A0(n537), .A1(readOutBus[334]), .B0(n536), .B1(
        readOutBus[454]), .Y(n522) );
  NAND4XLTS U911 ( .A(n525), .B(n524), .C(n523), .D(n522), .Y(readOut[34]) );
  AOI22X1TS U912 ( .A0(n531), .A1(readOutBus[33]), .B0(n530), .B1(
        readOutBus[153]), .Y(n529) );
  AOI22X1TS U913 ( .A0(n533), .A1(readOutBus[273]), .B0(n532), .B1(
        readOutBus[393]), .Y(n528) );
  AOI22X1TS U914 ( .A0(n535), .A1(readOutBus[93]), .B0(n534), .B1(
        readOutBus[213]), .Y(n527) );
  AOI22X1TS U915 ( .A0(n537), .A1(readOutBus[333]), .B0(n536), .B1(
        readOutBus[453]), .Y(n526) );
  NAND4XLTS U916 ( .A(n529), .B(n528), .C(n527), .D(n526), .Y(readOut[33]) );
  AOI22X1TS U917 ( .A0(n531), .A1(readOutBus[32]), .B0(n530), .B1(
        readOutBus[152]), .Y(n541) );
  AOI22X1TS U918 ( .A0(n533), .A1(readOutBus[272]), .B0(n532), .B1(
        readOutBus[392]), .Y(n540) );
  AOI22X1TS U919 ( .A0(n535), .A1(readOutBus[92]), .B0(n534), .B1(
        readOutBus[212]), .Y(n539) );
  AOI22X1TS U920 ( .A0(n537), .A1(readOutBus[332]), .B0(n536), .B1(
        readOutBus[452]), .Y(n538) );
  NAND4XLTS U921 ( .A(n541), .B(n540), .C(n539), .D(n538), .Y(readOut[32]) );
  CLKBUFX2TS U922 ( .A(n542), .Y(n559) );
  CLKBUFX2TS U923 ( .A(n586), .Y(n558) );
  AOI22X1TS U924 ( .A0(n559), .A1(readOutBus[31]), .B0(n558), .B1(
        readOutBus[151]), .Y(n549) );
  CLKBUFX2TS U925 ( .A(n543), .Y(n561) );
  CLKBUFX2TS U926 ( .A(n588), .Y(n560) );
  AOI22X1TS U927 ( .A0(n561), .A1(readOutBus[271]), .B0(n560), .B1(
        readOutBus[391]), .Y(n548) );
  CLKBUFX2TS U928 ( .A(n544), .Y(n563) );
  CLKBUFX2TS U929 ( .A(n590), .Y(n562) );
  AOI22X1TS U930 ( .A0(n563), .A1(readOutBus[91]), .B0(n562), .B1(
        readOutBus[211]), .Y(n547) );
  CLKBUFX2TS U931 ( .A(n545), .Y(n565) );
  CLKBUFX2TS U932 ( .A(n592), .Y(n564) );
  AOI22X1TS U933 ( .A0(n565), .A1(readOutBus[331]), .B0(n564), .B1(
        readOutBus[451]), .Y(n546) );
  NAND4XLTS U934 ( .A(n549), .B(n548), .C(n547), .D(n546), .Y(readOut[31]) );
  AOI22X1TS U935 ( .A0(n559), .A1(readOutBus[30]), .B0(n558), .B1(
        readOutBus[150]), .Y(n553) );
  AOI22X1TS U936 ( .A0(n561), .A1(readOutBus[270]), .B0(n560), .B1(
        readOutBus[390]), .Y(n552) );
  AOI22X1TS U937 ( .A0(n563), .A1(readOutBus[90]), .B0(n562), .B1(
        readOutBus[210]), .Y(n551) );
  AOI22X1TS U938 ( .A0(n565), .A1(readOutBus[330]), .B0(n564), .B1(
        readOutBus[450]), .Y(n550) );
  NAND4XLTS U939 ( .A(n553), .B(n552), .C(n551), .D(n550), .Y(readOut[30]) );
  AOI22X1TS U940 ( .A0(n559), .A1(readOutBus[29]), .B0(n558), .B1(
        readOutBus[149]), .Y(n557) );
  AOI22X1TS U941 ( .A0(n561), .A1(readOutBus[269]), .B0(n560), .B1(
        readOutBus[389]), .Y(n556) );
  AOI22X1TS U942 ( .A0(n563), .A1(readOutBus[89]), .B0(n562), .B1(
        readOutBus[209]), .Y(n555) );
  AOI22X1TS U943 ( .A0(n565), .A1(readOutBus[329]), .B0(n564), .B1(
        readOutBus[449]), .Y(n554) );
  NAND4XLTS U944 ( .A(n557), .B(n556), .C(n555), .D(n554), .Y(readOut[29]) );
  AOI22X1TS U945 ( .A0(n559), .A1(readOutBus[28]), .B0(n558), .B1(
        readOutBus[148]), .Y(n569) );
  AOI22X1TS U946 ( .A0(n561), .A1(readOutBus[268]), .B0(n560), .B1(
        readOutBus[388]), .Y(n568) );
  AOI22X1TS U947 ( .A0(n563), .A1(readOutBus[88]), .B0(n562), .B1(
        readOutBus[208]), .Y(n567) );
  AOI22X1TS U948 ( .A0(n565), .A1(readOutBus[328]), .B0(n564), .B1(
        readOutBus[448]), .Y(n566) );
  NAND4XLTS U949 ( .A(n569), .B(n568), .C(n567), .D(n566), .Y(readOut[28]) );
  CLKBUFX2TS U950 ( .A(n626), .Y(n587) );
  AOI22X1TS U951 ( .A0(n587), .A1(readOutBus[27]), .B0(n627), .B1(
        readOutBus[147]), .Y(n573) );
  CLKBUFX2TS U952 ( .A(n628), .Y(n589) );
  AOI22X1TS U953 ( .A0(n589), .A1(readOutBus[267]), .B0(n629), .B1(
        readOutBus[387]), .Y(n572) );
  CLKBUFX2TS U954 ( .A(n630), .Y(n591) );
  AOI22X1TS U955 ( .A0(n591), .A1(readOutBus[87]), .B0(n631), .B1(
        readOutBus[207]), .Y(n571) );
  CLKBUFX2TS U956 ( .A(n632), .Y(n593) );
  AOI22X1TS U957 ( .A0(n593), .A1(readOutBus[327]), .B0(n633), .B1(
        readOutBus[447]), .Y(n570) );
  NAND4XLTS U958 ( .A(n573), .B(n572), .C(n571), .D(n570), .Y(readOut[27]) );
  CLKBUFX2TS U959 ( .A(n598), .Y(n735) );
  AOI22X1TS U960 ( .A0(n587), .A1(readOutBus[26]), .B0(n735), .B1(
        readOutBus[146]), .Y(n577) );
  CLKBUFX2TS U961 ( .A(n599), .Y(n737) );
  AOI22X1TS U962 ( .A0(n589), .A1(readOutBus[266]), .B0(n737), .B1(
        readOutBus[386]), .Y(n576) );
  CLKBUFX2TS U963 ( .A(n631), .Y(n739) );
  AOI22X1TS U964 ( .A0(n591), .A1(readOutBus[86]), .B0(n739), .B1(
        readOutBus[206]), .Y(n575) );
  CLKBUFX2TS U965 ( .A(n601), .Y(n741) );
  AOI22X1TS U966 ( .A0(n593), .A1(readOutBus[326]), .B0(n741), .B1(
        readOutBus[446]), .Y(n574) );
  NAND4XLTS U967 ( .A(n577), .B(n576), .C(n575), .D(n574), .Y(readOut[26]) );
  AOI22X1TS U968 ( .A0(n587), .A1(readOutBus[25]), .B0(n578), .B1(
        readOutBus[145]), .Y(n585) );
  AOI22X1TS U969 ( .A0(n589), .A1(readOutBus[265]), .B0(n579), .B1(
        readOutBus[385]), .Y(n584) );
  AOI22X1TS U970 ( .A0(n591), .A1(readOutBus[85]), .B0(n580), .B1(
        readOutBus[205]), .Y(n583) );
  AOI22X1TS U971 ( .A0(n593), .A1(readOutBus[325]), .B0(n581), .B1(
        readOutBus[445]), .Y(n582) );
  NAND4XLTS U972 ( .A(n585), .B(n584), .C(n583), .D(n582), .Y(readOut[25]) );
  AOI22X1TS U973 ( .A0(n587), .A1(readOutBus[24]), .B0(n586), .B1(
        readOutBus[144]), .Y(n597) );
  AOI22X1TS U974 ( .A0(n589), .A1(readOutBus[264]), .B0(n588), .B1(
        readOutBus[384]), .Y(n596) );
  AOI22X1TS U975 ( .A0(n591), .A1(readOutBus[84]), .B0(n590), .B1(
        readOutBus[204]), .Y(n595) );
  AOI22X1TS U976 ( .A0(n593), .A1(readOutBus[324]), .B0(n592), .B1(
        readOutBus[444]), .Y(n594) );
  NAND4XLTS U977 ( .A(n597), .B(n596), .C(n595), .D(n594), .Y(readOut[24]) );
  CLKBUFX2TS U978 ( .A(n734), .Y(n615) );
  CLKBUFX2TS U979 ( .A(n598), .Y(n614) );
  AOI22X1TS U980 ( .A0(n615), .A1(readOutBus[23]), .B0(n614), .B1(
        readOutBus[143]), .Y(n605) );
  CLKBUFX2TS U981 ( .A(n736), .Y(n617) );
  CLKBUFX2TS U982 ( .A(n599), .Y(n616) );
  AOI22X1TS U983 ( .A0(n617), .A1(readOutBus[263]), .B0(n616), .B1(
        readOutBus[383]), .Y(n604) );
  CLKBUFX2TS U984 ( .A(n738), .Y(n619) );
  CLKBUFX2TS U985 ( .A(n600), .Y(n618) );
  AOI22X1TS U986 ( .A0(n619), .A1(readOutBus[83]), .B0(n618), .B1(
        readOutBus[203]), .Y(n603) );
  CLKBUFX2TS U987 ( .A(n740), .Y(n621) );
  CLKBUFX2TS U988 ( .A(n601), .Y(n620) );
  AOI22X1TS U989 ( .A0(n621), .A1(readOutBus[323]), .B0(n620), .B1(
        readOutBus[443]), .Y(n602) );
  NAND4XLTS U990 ( .A(n605), .B(n604), .C(n603), .D(n602), .Y(readOut[23]) );
  AOI22X1TS U991 ( .A0(n615), .A1(readOutBus[22]), .B0(n614), .B1(
        readOutBus[142]), .Y(n609) );
  AOI22X1TS U992 ( .A0(n617), .A1(readOutBus[262]), .B0(n616), .B1(
        readOutBus[382]), .Y(n608) );
  AOI22X1TS U993 ( .A0(n619), .A1(readOutBus[82]), .B0(n618), .B1(
        readOutBus[202]), .Y(n607) );
  AOI22X1TS U994 ( .A0(n621), .A1(readOutBus[322]), .B0(n620), .B1(
        readOutBus[442]), .Y(n606) );
  NAND4XLTS U995 ( .A(n609), .B(n608), .C(n607), .D(n606), .Y(readOut[22]) );
  AOI22X1TS U996 ( .A0(n615), .A1(readOutBus[21]), .B0(n614), .B1(
        readOutBus[141]), .Y(n613) );
  AOI22X1TS U997 ( .A0(n617), .A1(readOutBus[261]), .B0(n616), .B1(
        readOutBus[381]), .Y(n612) );
  AOI22X1TS U998 ( .A0(n619), .A1(readOutBus[81]), .B0(n618), .B1(
        readOutBus[201]), .Y(n611) );
  AOI22X1TS U999 ( .A0(n621), .A1(readOutBus[321]), .B0(n620), .B1(
        readOutBus[441]), .Y(n610) );
  NAND4XLTS U1000 ( .A(n613), .B(n612), .C(n611), .D(n610), .Y(readOut[21]) );
  AOI22X1TS U1001 ( .A0(n615), .A1(readOutBus[20]), .B0(n614), .B1(
        readOutBus[140]), .Y(n625) );
  AOI22X1TS U1002 ( .A0(n617), .A1(readOutBus[260]), .B0(n616), .B1(
        readOutBus[380]), .Y(n624) );
  AOI22X1TS U1003 ( .A0(n619), .A1(readOutBus[80]), .B0(n618), .B1(
        readOutBus[200]), .Y(n623) );
  AOI22X1TS U1004 ( .A0(n621), .A1(readOutBus[320]), .B0(n620), .B1(
        readOutBus[440]), .Y(n622) );
  NAND4XLTS U1005 ( .A(n625), .B(n624), .C(n623), .D(n622), .Y(readOut[20]) );
  CLKBUFX2TS U1006 ( .A(n626), .Y(n647) );
  CLKBUFX2TS U1007 ( .A(n627), .Y(n646) );
  AOI22X1TS U1008 ( .A0(n647), .A1(readOutBus[19]), .B0(n646), .B1(
        readOutBus[139]), .Y(n637) );
  CLKBUFX2TS U1009 ( .A(n628), .Y(n649) );
  CLKBUFX2TS U1010 ( .A(n629), .Y(n648) );
  AOI22X1TS U1011 ( .A0(n649), .A1(readOutBus[259]), .B0(n648), .B1(
        readOutBus[379]), .Y(n636) );
  CLKBUFX2TS U1012 ( .A(n630), .Y(n651) );
  CLKBUFX2TS U1013 ( .A(n631), .Y(n650) );
  AOI22X1TS U1014 ( .A0(n651), .A1(readOutBus[79]), .B0(n650), .B1(
        readOutBus[199]), .Y(n635) );
  CLKBUFX2TS U1015 ( .A(n632), .Y(n653) );
  CLKBUFX2TS U1016 ( .A(n633), .Y(n652) );
  AOI22X1TS U1017 ( .A0(n653), .A1(readOutBus[319]), .B0(n652), .B1(
        readOutBus[439]), .Y(n634) );
  NAND4XLTS U1018 ( .A(n637), .B(n636), .C(n635), .D(n634), .Y(readOut[19]) );
  AOI22X1TS U1019 ( .A0(n647), .A1(readOutBus[18]), .B0(n646), .B1(
        readOutBus[138]), .Y(n641) );
  AOI22X1TS U1020 ( .A0(n649), .A1(readOutBus[258]), .B0(n648), .B1(
        readOutBus[378]), .Y(n640) );
  AOI22X1TS U1021 ( .A0(n651), .A1(readOutBus[78]), .B0(n650), .B1(
        readOutBus[198]), .Y(n639) );
  AOI22X1TS U1022 ( .A0(n653), .A1(readOutBus[318]), .B0(n652), .B1(
        readOutBus[438]), .Y(n638) );
  NAND4XLTS U1023 ( .A(n641), .B(n640), .C(n639), .D(n638), .Y(readOut[18]) );
  AOI22X1TS U1024 ( .A0(n647), .A1(readOutBus[17]), .B0(n646), .B1(
        readOutBus[137]), .Y(n645) );
  AOI22X1TS U1025 ( .A0(n649), .A1(readOutBus[257]), .B0(n648), .B1(
        readOutBus[377]), .Y(n644) );
  AOI22X1TS U1026 ( .A0(n651), .A1(readOutBus[77]), .B0(n650), .B1(
        readOutBus[197]), .Y(n643) );
  AOI22X1TS U1027 ( .A0(n653), .A1(readOutBus[317]), .B0(n652), .B1(
        readOutBus[437]), .Y(n642) );
  NAND4XLTS U1028 ( .A(n645), .B(n644), .C(n643), .D(n642), .Y(readOut[17]) );
  AOI22X1TS U1029 ( .A0(n647), .A1(readOutBus[16]), .B0(n646), .B1(
        readOutBus[136]), .Y(n657) );
  AOI22X1TS U1030 ( .A0(n649), .A1(readOutBus[256]), .B0(n648), .B1(
        readOutBus[376]), .Y(n656) );
  AOI22X1TS U1031 ( .A0(n651), .A1(readOutBus[76]), .B0(n650), .B1(
        readOutBus[196]), .Y(n655) );
  AOI22X1TS U1032 ( .A0(n653), .A1(readOutBus[316]), .B0(n652), .B1(
        readOutBus[436]), .Y(n654) );
  NAND4XLTS U1033 ( .A(n657), .B(n656), .C(n655), .D(n654), .Y(readOut[16]) );
  CLKBUFX2TS U1034 ( .A(n706), .Y(n671) );
  CLKBUFX2TS U1035 ( .A(n735), .Y(n670) );
  AOI22X1TS U1036 ( .A0(n671), .A1(readOutBus[15]), .B0(n670), .B1(
        readOutBus[135]), .Y(n661) );
  CLKBUFX2TS U1037 ( .A(n708), .Y(n673) );
  CLKBUFX2TS U1038 ( .A(n737), .Y(n672) );
  AOI22X1TS U1039 ( .A0(n673), .A1(readOutBus[255]), .B0(n672), .B1(
        readOutBus[375]), .Y(n660) );
  CLKBUFX2TS U1040 ( .A(n710), .Y(n675) );
  CLKBUFX2TS U1041 ( .A(n739), .Y(n674) );
  AOI22X1TS U1042 ( .A0(n675), .A1(readOutBus[75]), .B0(n674), .B1(
        readOutBus[195]), .Y(n659) );
  CLKBUFX2TS U1043 ( .A(n712), .Y(n677) );
  CLKBUFX2TS U1044 ( .A(n741), .Y(n676) );
  AOI22X1TS U1045 ( .A0(n677), .A1(readOutBus[315]), .B0(n676), .B1(
        readOutBus[435]), .Y(n658) );
  NAND4XLTS U1046 ( .A(n661), .B(n660), .C(n659), .D(n658), .Y(readOut[15]) );
  AOI22X1TS U1047 ( .A0(n671), .A1(readOutBus[14]), .B0(n670), .B1(
        readOutBus[134]), .Y(n665) );
  AOI22X1TS U1048 ( .A0(n673), .A1(readOutBus[254]), .B0(n672), .B1(
        readOutBus[374]), .Y(n664) );
  AOI22X1TS U1049 ( .A0(n675), .A1(readOutBus[74]), .B0(n674), .B1(
        readOutBus[194]), .Y(n663) );
  AOI22X1TS U1050 ( .A0(n677), .A1(readOutBus[314]), .B0(n676), .B1(
        readOutBus[434]), .Y(n662) );
  NAND4XLTS U1051 ( .A(n665), .B(n664), .C(n663), .D(n662), .Y(readOut[14]) );
  AOI22X1TS U1052 ( .A0(n671), .A1(readOutBus[13]), .B0(n670), .B1(
        readOutBus[133]), .Y(n669) );
  AOI22X1TS U1053 ( .A0(n673), .A1(readOutBus[253]), .B0(n672), .B1(
        readOutBus[373]), .Y(n668) );
  AOI22X1TS U1054 ( .A0(n675), .A1(readOutBus[73]), .B0(n674), .B1(
        readOutBus[193]), .Y(n667) );
  AOI22X1TS U1055 ( .A0(n677), .A1(readOutBus[313]), .B0(n676), .B1(
        readOutBus[433]), .Y(n666) );
  NAND4XLTS U1056 ( .A(n669), .B(n668), .C(n667), .D(n666), .Y(readOut[13]) );
  AOI22X1TS U1057 ( .A0(n671), .A1(readOutBus[12]), .B0(n670), .B1(
        readOutBus[132]), .Y(n681) );
  AOI22X1TS U1058 ( .A0(n673), .A1(readOutBus[252]), .B0(n672), .B1(
        readOutBus[372]), .Y(n680) );
  AOI22X1TS U1059 ( .A0(n675), .A1(readOutBus[72]), .B0(n674), .B1(
        readOutBus[192]), .Y(n679) );
  AOI22X1TS U1060 ( .A0(n677), .A1(readOutBus[312]), .B0(n676), .B1(
        readOutBus[432]), .Y(n678) );
  NAND4XLTS U1061 ( .A(n681), .B(n680), .C(n679), .D(n678), .Y(readOut[12]) );
  CLKBUFX2TS U1062 ( .A(n706), .Y(n695) );
  CLKBUFX2TS U1063 ( .A(n735), .Y(n694) );
  AOI22X1TS U1064 ( .A0(n695), .A1(readOutBus[11]), .B0(n694), .B1(
        readOutBus[131]), .Y(n685) );
  CLKBUFX2TS U1065 ( .A(n708), .Y(n697) );
  CLKBUFX2TS U1066 ( .A(n737), .Y(n696) );
  AOI22X1TS U1067 ( .A0(n697), .A1(readOutBus[251]), .B0(n696), .B1(
        readOutBus[371]), .Y(n684) );
  CLKBUFX2TS U1068 ( .A(n710), .Y(n699) );
  CLKBUFX2TS U1069 ( .A(n739), .Y(n698) );
  AOI22X1TS U1070 ( .A0(n699), .A1(readOutBus[71]), .B0(n698), .B1(
        readOutBus[191]), .Y(n683) );
  CLKBUFX2TS U1071 ( .A(n712), .Y(n701) );
  CLKBUFX2TS U1072 ( .A(n741), .Y(n700) );
  AOI22X1TS U1073 ( .A0(n701), .A1(readOutBus[311]), .B0(n700), .B1(
        readOutBus[431]), .Y(n682) );
  NAND4XLTS U1074 ( .A(n685), .B(n684), .C(n683), .D(n682), .Y(readOut[11]) );
  AOI22X1TS U1075 ( .A0(n695), .A1(readOutBus[10]), .B0(n694), .B1(
        readOutBus[130]), .Y(n689) );
  AOI22X1TS U1076 ( .A0(n697), .A1(readOutBus[250]), .B0(n696), .B1(
        readOutBus[370]), .Y(n688) );
  AOI22X1TS U1077 ( .A0(n699), .A1(readOutBus[70]), .B0(n698), .B1(
        readOutBus[190]), .Y(n687) );
  AOI22X1TS U1078 ( .A0(n701), .A1(readOutBus[310]), .B0(n700), .B1(
        readOutBus[430]), .Y(n686) );
  NAND4XLTS U1079 ( .A(n689), .B(n688), .C(n687), .D(n686), .Y(readOut[10]) );
  AOI22X1TS U1080 ( .A0(n695), .A1(readOutBus[9]), .B0(n694), .B1(
        readOutBus[129]), .Y(n693) );
  AOI22X1TS U1081 ( .A0(n697), .A1(readOutBus[249]), .B0(n696), .B1(
        readOutBus[369]), .Y(n692) );
  AOI22X1TS U1082 ( .A0(n699), .A1(readOutBus[69]), .B0(n698), .B1(
        readOutBus[189]), .Y(n691) );
  AOI22X1TS U1083 ( .A0(n701), .A1(readOutBus[309]), .B0(n700), .B1(
        readOutBus[429]), .Y(n690) );
  NAND4XLTS U1084 ( .A(n693), .B(n692), .C(n691), .D(n690), .Y(readOut[9]) );
  AOI22X1TS U1085 ( .A0(n695), .A1(readOutBus[8]), .B0(n694), .B1(
        readOutBus[128]), .Y(n705) );
  AOI22X1TS U1086 ( .A0(n697), .A1(readOutBus[248]), .B0(n696), .B1(
        readOutBus[368]), .Y(n704) );
  AOI22X1TS U1087 ( .A0(n699), .A1(readOutBus[68]), .B0(n698), .B1(
        readOutBus[188]), .Y(n703) );
  AOI22X1TS U1088 ( .A0(n701), .A1(readOutBus[308]), .B0(n700), .B1(
        readOutBus[428]), .Y(n702) );
  NAND4XLTS U1089 ( .A(n705), .B(n704), .C(n703), .D(n702), .Y(readOut[8]) );
  CLKBUFX2TS U1090 ( .A(n707), .Y(n726) );
  AOI22X1TS U1091 ( .A0(n414), .A1(readOutBus[7]), .B0(n726), .B1(
        readOutBus[127]), .Y(n717) );
  CLKBUFX2TS U1092 ( .A(n709), .Y(n727) );
  AOI22X1TS U1093 ( .A0(n415), .A1(readOutBus[247]), .B0(n727), .B1(
        readOutBus[367]), .Y(n716) );
  CLKBUFX2TS U1094 ( .A(n711), .Y(n728) );
  AOI22X1TS U1095 ( .A0(n416), .A1(readOutBus[67]), .B0(n728), .B1(
        readOutBus[187]), .Y(n715) );
  CLKBUFX2TS U1096 ( .A(n713), .Y(n729) );
  AOI22X1TS U1097 ( .A0(n417), .A1(readOutBus[307]), .B0(n729), .B1(
        readOutBus[427]), .Y(n714) );
  NAND4XLTS U1098 ( .A(n717), .B(n716), .C(n715), .D(n714), .Y(readOut[7]) );
  AOI22X1TS U1099 ( .A0(n542), .A1(readOutBus[6]), .B0(n726), .B1(
        readOutBus[126]), .Y(n721) );
  AOI22X1TS U1100 ( .A0(n543), .A1(readOutBus[246]), .B0(n727), .B1(
        readOutBus[366]), .Y(n720) );
  AOI22X1TS U1101 ( .A0(n544), .A1(readOutBus[66]), .B0(n728), .B1(
        readOutBus[186]), .Y(n719) );
  AOI22X1TS U1102 ( .A0(n545), .A1(readOutBus[306]), .B0(n729), .B1(
        readOutBus[426]), .Y(n718) );
  NAND4XLTS U1103 ( .A(n721), .B(n720), .C(n719), .D(n718), .Y(readOut[6]) );
  AOI22X1TS U1104 ( .A0(n706), .A1(readOutBus[5]), .B0(n726), .B1(
        readOutBus[125]), .Y(n725) );
  AOI22X1TS U1105 ( .A0(n708), .A1(readOutBus[245]), .B0(n727), .B1(
        readOutBus[365]), .Y(n724) );
  AOI22X1TS U1106 ( .A0(n710), .A1(readOutBus[65]), .B0(n728), .B1(
        readOutBus[185]), .Y(n723) );
  AOI22X1TS U1107 ( .A0(n712), .A1(readOutBus[305]), .B0(n729), .B1(
        readOutBus[425]), .Y(n722) );
  NAND4XLTS U1108 ( .A(n725), .B(n724), .C(n723), .D(n722), .Y(readOut[5]) );
  AOI22X1TS U1109 ( .A0(n414), .A1(readOutBus[4]), .B0(n726), .B1(
        readOutBus[124]), .Y(n733) );
  AOI22X1TS U1110 ( .A0(n415), .A1(readOutBus[244]), .B0(n727), .B1(
        readOutBus[364]), .Y(n732) );
  AOI22X1TS U1111 ( .A0(n416), .A1(readOutBus[64]), .B0(n728), .B1(
        readOutBus[184]), .Y(n731) );
  AOI22X1TS U1112 ( .A0(n417), .A1(readOutBus[304]), .B0(n729), .B1(
        readOutBus[424]), .Y(n730) );
  NAND4XLTS U1113 ( .A(n733), .B(n732), .C(n731), .D(n730), .Y(readOut[4]) );
  CLKBUFX2TS U1114 ( .A(n734), .Y(n755) );
  CLKBUFX2TS U1115 ( .A(n735), .Y(n754) );
  AOI22X1TS U1116 ( .A0(n755), .A1(readOutBus[3]), .B0(n754), .B1(
        readOutBus[123]), .Y(n745) );
  CLKBUFX2TS U1117 ( .A(n736), .Y(n757) );
  CLKBUFX2TS U1118 ( .A(n737), .Y(n756) );
  AOI22X1TS U1119 ( .A0(n757), .A1(readOutBus[243]), .B0(n756), .B1(
        readOutBus[363]), .Y(n744) );
  CLKBUFX2TS U1120 ( .A(n738), .Y(n759) );
  CLKBUFX2TS U1121 ( .A(n739), .Y(n758) );
  AOI22X1TS U1122 ( .A0(n759), .A1(readOutBus[63]), .B0(n758), .B1(
        readOutBus[183]), .Y(n743) );
  CLKBUFX2TS U1123 ( .A(n740), .Y(n761) );
  CLKBUFX2TS U1124 ( .A(n741), .Y(n760) );
  AOI22X1TS U1125 ( .A0(n761), .A1(readOutBus[303]), .B0(n760), .B1(
        readOutBus[423]), .Y(n742) );
  NAND4XLTS U1126 ( .A(n745), .B(n744), .C(n743), .D(n742), .Y(readOut[3]) );
  AOI22X1TS U1127 ( .A0(n755), .A1(readOutBus[2]), .B0(n754), .B1(
        readOutBus[122]), .Y(n749) );
  AOI22X1TS U1128 ( .A0(n757), .A1(readOutBus[242]), .B0(n756), .B1(
        readOutBus[362]), .Y(n748) );
  AOI22X1TS U1129 ( .A0(n759), .A1(readOutBus[62]), .B0(n758), .B1(
        readOutBus[182]), .Y(n747) );
  AOI22X1TS U1130 ( .A0(n761), .A1(readOutBus[302]), .B0(n760), .B1(
        readOutBus[422]), .Y(n746) );
  NAND4XLTS U1131 ( .A(n749), .B(n748), .C(n747), .D(n746), .Y(readOut[2]) );
  AOI22X1TS U1132 ( .A0(n755), .A1(readOutBus[1]), .B0(n754), .B1(
        readOutBus[121]), .Y(n753) );
  AOI22X1TS U1133 ( .A0(n757), .A1(readOutBus[241]), .B0(n756), .B1(
        readOutBus[361]), .Y(n752) );
  AOI22X1TS U1134 ( .A0(n759), .A1(readOutBus[61]), .B0(n758), .B1(
        readOutBus[181]), .Y(n751) );
  AOI22X1TS U1135 ( .A0(n761), .A1(readOutBus[301]), .B0(n760), .B1(
        readOutBus[421]), .Y(n750) );
  NAND4XLTS U1136 ( .A(n753), .B(n752), .C(n751), .D(n750), .Y(readOut[1]) );
  AOI22X1TS U1137 ( .A0(n755), .A1(readOutBus[0]), .B0(n754), .B1(
        readOutBus[120]), .Y(n765) );
  AOI22X1TS U1138 ( .A0(n757), .A1(readOutBus[240]), .B0(n756), .B1(
        readOutBus[360]), .Y(n764) );
  AOI22X1TS U1139 ( .A0(n759), .A1(readOutBus[60]), .B0(n758), .B1(
        readOutBus[180]), .Y(n763) );
  AOI22X1TS U1140 ( .A0(n761), .A1(readOutBus[300]), .B0(n760), .B1(
        readOutBus[420]), .Y(n762) );
  NAND4XLTS U1141 ( .A(n765), .B(n764), .C(n763), .D(n762), .Y(readOut[0]) );
endmodule

