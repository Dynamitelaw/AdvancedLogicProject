
module Layer1WeightStorage ( writeEnable, NodeSelect, writeIn, readOut );
  input [9:0] NodeSelect;
  input [159:0] writeIn;
  output [159:0] readOut;
  input writeEnable;
  wire   n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107;
  wire   [959:0] readOutBus;

  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_44_ ( .G(n1907), .D(n1637), 
        .Q(readOutBus[44]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_45_ ( .G(n1907), .D(n1639), 
        .Q(readOutBus[45]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_46_ ( .G(n1907), .D(n1641), 
        .Q(readOutBus[46]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_47_ ( .G(n1907), .D(n1643), 
        .Q(readOutBus[47]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_76_ ( .G(n1899), .D(n1701), 
        .Q(readOutBus[76]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_77_ ( .G(n1899), .D(n1703), 
        .Q(readOutBus[77]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_78_ ( .G(n1899), .D(n1705), 
        .Q(readOutBus[78]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_79_ ( .G(n1899), .D(n1707), 
        .Q(readOutBus[79]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_84_ ( .G(n1897), .D(n1717), 
        .Q(readOutBus[84]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_85_ ( .G(n1897), .D(n1719), 
        .Q(readOutBus[85]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_86_ ( .G(n1897), .D(n1721), 
        .Q(readOutBus[86]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_87_ ( .G(n1897), .D(n1723), 
        .Q(readOutBus[87]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_88_ ( .G(n1896), .D(n1725), 
        .Q(readOutBus[88]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_89_ ( .G(n1896), .D(n1727), 
        .Q(readOutBus[89]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_90_ ( .G(n1896), .D(n1729), 
        .Q(readOutBus[90]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_91_ ( .G(n1896), .D(n1731), 
        .Q(readOutBus[91]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_92_ ( .G(n1895), .D(n1733), 
        .Q(readOutBus[92]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_93_ ( .G(n1895), .D(n1735), 
        .Q(readOutBus[93]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_94_ ( .G(n1895), .D(n1737), 
        .Q(readOutBus[94]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_95_ ( .G(n1895), .D(n1739), 
        .Q(readOutBus[95]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_120_ ( .G(n722), .D(n1789), 
        .Q(readOutBus[120]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_121_ ( .G(n723), .D(n1791), 
        .Q(readOutBus[121]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_122_ ( .G(n706), .D(n1793), 
        .Q(readOutBus[122]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_123_ ( .G(n707), .D(n1795), 
        .Q(readOutBus[123]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_124_ ( .G(n1888), .D(n1797), 
        .Q(readOutBus[124]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_125_ ( .G(n1888), .D(n1799), 
        .Q(readOutBus[125]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_126_ ( .G(n1888), .D(n1801), 
        .Q(readOutBus[126]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_127_ ( .G(n1888), .D(n1803), 
        .Q(readOutBus[127]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_128_ ( .G(n1887), .D(n1805), 
        .Q(readOutBus[128]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_129_ ( .G(n1887), .D(n1807), 
        .Q(readOutBus[129]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_130_ ( .G(n1887), .D(n1809), 
        .Q(readOutBus[130]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_131_ ( .G(n1887), .D(n1811), 
        .Q(readOutBus[131]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_132_ ( .G(n1886), .D(n1813), 
        .Q(readOutBus[132]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_133_ ( .G(n1886), .D(n1815), 
        .Q(readOutBus[133]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_134_ ( .G(n1886), .D(n1817), 
        .Q(readOutBus[134]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_135_ ( .G(n1886), .D(n1819), 
        .Q(readOutBus[135]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_136_ ( .G(n1885), .D(n1821), 
        .Q(readOutBus[136]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_137_ ( .G(n1885), .D(n1823), 
        .Q(readOutBus[137]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_138_ ( .G(n1885), .D(n1825), 
        .Q(readOutBus[138]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_139_ ( .G(n1885), .D(n1827), 
        .Q(readOutBus[139]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_140_ ( .G(n1884), .D(n1829), 
        .Q(readOutBus[140]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_141_ ( .G(n1884), .D(n1831), 
        .Q(readOutBus[141]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_142_ ( .G(n1884), .D(n1833), 
        .Q(readOutBus[142]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_143_ ( .G(n1884), .D(n1835), 
        .Q(readOutBus[143]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_144_ ( .G(n1883), .D(n1837), 
        .Q(readOutBus[144]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_145_ ( .G(n1883), .D(n1839), 
        .Q(readOutBus[145]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_146_ ( .G(n1883), .D(n1841), 
        .Q(readOutBus[146]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_147_ ( .G(n1883), .D(n1843), 
        .Q(readOutBus[147]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_152_ ( .G(n1881), .D(n1853), 
        .Q(readOutBus[152]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_153_ ( .G(n1881), .D(n1855), 
        .Q(readOutBus[153]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_154_ ( .G(n1881), .D(n1857), 
        .Q(readOutBus[154]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_155_ ( .G(n1881), .D(n1859), 
        .Q(readOutBus[155]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_156_ ( .G(n1880), .D(n1861), 
        .Q(readOutBus[156]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_157_ ( .G(n1880), .D(n1863), 
        .Q(readOutBus[157]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_158_ ( .G(n1880), .D(n1865), 
        .Q(readOutBus[158]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_159_ ( .G(n1880), .D(n1867), 
        .Q(readOutBus[159]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_44_ ( .G(n1983), .D(n1637), 
        .Q(readOutBus[364]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_45_ ( .G(n1983), .D(n1639), 
        .Q(readOutBus[365]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_46_ ( .G(n1983), .D(n1641), 
        .Q(readOutBus[366]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_47_ ( .G(n1983), .D(n1643), 
        .Q(readOutBus[367]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_76_ ( .G(n1975), .D(n1701), 
        .Q(readOutBus[396]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_77_ ( .G(n1975), .D(n1703), 
        .Q(readOutBus[397]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_78_ ( .G(n1975), .D(n1705), 
        .Q(readOutBus[398]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_79_ ( .G(n1975), .D(n1707), 
        .Q(readOutBus[399]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_84_ ( .G(n1973), .D(n1717), 
        .Q(readOutBus[404]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_85_ ( .G(n1973), .D(n1719), 
        .Q(readOutBus[405]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_86_ ( .G(n1973), .D(n1721), 
        .Q(readOutBus[406]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_87_ ( .G(n1973), .D(n1723), 
        .Q(readOutBus[407]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_88_ ( .G(n1972), .D(n1725), 
        .Q(readOutBus[408]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_89_ ( .G(n1972), .D(n1727), 
        .Q(readOutBus[409]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_90_ ( .G(n1972), .D(n1729), 
        .Q(readOutBus[410]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_91_ ( .G(n1972), .D(n1731), 
        .Q(readOutBus[411]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_92_ ( .G(n1971), .D(n1733), 
        .Q(readOutBus[412]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_93_ ( .G(n1971), .D(n1735), 
        .Q(readOutBus[413]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_94_ ( .G(n1971), .D(n1737), 
        .Q(readOutBus[414]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_95_ ( .G(n1971), .D(n1739), 
        .Q(readOutBus[415]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_120_ ( .G(n720), .D(n1789), 
        .Q(readOutBus[440]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_121_ ( .G(n721), .D(n1791), 
        .Q(readOutBus[441]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_122_ ( .G(n704), .D(n1793), 
        .Q(readOutBus[442]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_123_ ( .G(n705), .D(n1795), 
        .Q(readOutBus[443]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_124_ ( .G(n1964), .D(n1797), 
        .Q(readOutBus[444]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_125_ ( .G(n1964), .D(n1799), 
        .Q(readOutBus[445]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_126_ ( .G(n1964), .D(n1801), 
        .Q(readOutBus[446]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_127_ ( .G(n1964), .D(n1803), 
        .Q(readOutBus[447]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_128_ ( .G(n1963), .D(n1805), 
        .Q(readOutBus[448]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_129_ ( .G(n1963), .D(n1807), 
        .Q(readOutBus[449]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_130_ ( .G(n1963), .D(n1809), 
        .Q(readOutBus[450]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_131_ ( .G(n1963), .D(n1811), 
        .Q(readOutBus[451]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_132_ ( .G(n1962), .D(n1813), 
        .Q(readOutBus[452]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_133_ ( .G(n1962), .D(n1815), 
        .Q(readOutBus[453]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_134_ ( .G(n1962), .D(n1817), 
        .Q(readOutBus[454]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_135_ ( .G(n1962), .D(n1819), 
        .Q(readOutBus[455]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_136_ ( .G(n1961), .D(n1821), 
        .Q(readOutBus[456]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_137_ ( .G(n1961), .D(n1823), 
        .Q(readOutBus[457]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_138_ ( .G(n1961), .D(n1825), 
        .Q(readOutBus[458]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_139_ ( .G(n1961), .D(n1827), 
        .Q(readOutBus[459]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_140_ ( .G(n1960), .D(n1829), 
        .Q(readOutBus[460]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_141_ ( .G(n1960), .D(n1831), 
        .Q(readOutBus[461]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_142_ ( .G(n1960), .D(n1833), 
        .Q(readOutBus[462]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_143_ ( .G(n1960), .D(n1835), 
        .Q(readOutBus[463]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_144_ ( .G(n1959), .D(n1837), 
        .Q(readOutBus[464]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_145_ ( .G(n1959), .D(n1839), 
        .Q(readOutBus[465]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_146_ ( .G(n1959), .D(n1841), 
        .Q(readOutBus[466]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_147_ ( .G(n1959), .D(n1843), 
        .Q(readOutBus[467]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_152_ ( .G(n1957), .D(n1853), 
        .Q(readOutBus[472]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_153_ ( .G(n1957), .D(n1855), 
        .Q(readOutBus[473]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_154_ ( .G(n1957), .D(n1857), 
        .Q(readOutBus[474]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_155_ ( .G(n1957), .D(n1859), 
        .Q(readOutBus[475]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_156_ ( .G(n1956), .D(n1861), 
        .Q(readOutBus[476]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_157_ ( .G(n1956), .D(n1863), 
        .Q(readOutBus[477]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_158_ ( .G(n1956), .D(n1865), 
        .Q(readOutBus[478]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_159_ ( .G(n1956), .D(n1867), 
        .Q(readOutBus[479]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_44_ ( .G(n2059), .D(n1637), 
        .Q(readOutBus[684]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_45_ ( .G(n2059), .D(n1639), 
        .Q(readOutBus[685]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_46_ ( .G(n2059), .D(n1641), 
        .Q(readOutBus[686]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_47_ ( .G(n2059), .D(n1643), 
        .Q(readOutBus[687]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_76_ ( .G(n2051), .D(n1701), 
        .Q(readOutBus[716]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_77_ ( .G(n2051), .D(n1703), 
        .Q(readOutBus[717]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_78_ ( .G(n2051), .D(n1705), 
        .Q(readOutBus[718]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_79_ ( .G(n2051), .D(n1707), 
        .Q(readOutBus[719]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_84_ ( .G(n2049), .D(n1717), 
        .Q(readOutBus[724]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_85_ ( .G(n2049), .D(n1719), 
        .Q(readOutBus[725]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_86_ ( .G(n2049), .D(n1721), 
        .Q(readOutBus[726]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_87_ ( .G(n2049), .D(n1723), 
        .Q(readOutBus[727]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_88_ ( .G(n2048), .D(n1725), 
        .Q(readOutBus[728]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_89_ ( .G(n2048), .D(n1727), 
        .Q(readOutBus[729]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_90_ ( .G(n2048), .D(n1729), 
        .Q(readOutBus[730]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_91_ ( .G(n2048), .D(n1731), 
        .Q(readOutBus[731]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_92_ ( .G(n2047), .D(n1733), 
        .Q(readOutBus[732]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_93_ ( .G(n2047), .D(n1735), 
        .Q(readOutBus[733]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_94_ ( .G(n2047), .D(n1737), 
        .Q(readOutBus[734]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_95_ ( .G(n2047), .D(n1739), 
        .Q(readOutBus[735]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_120_ ( .G(n724), .D(n1789), 
        .Q(readOutBus[760]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_121_ ( .G(n698), .D(n1791), 
        .Q(readOutBus[761]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_122_ ( .G(n710), .D(n1793), 
        .Q(readOutBus[762]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_123_ ( .G(n711), .D(n1795), 
        .Q(readOutBus[763]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_124_ ( .G(n2040), .D(n1797), 
        .Q(readOutBus[764]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_125_ ( .G(n2040), .D(n1799), 
        .Q(readOutBus[765]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_126_ ( .G(n2040), .D(n1801), 
        .Q(readOutBus[766]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_127_ ( .G(n2040), .D(n1803), 
        .Q(readOutBus[767]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_128_ ( .G(n2039), .D(n1805), 
        .Q(readOutBus[768]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_129_ ( .G(n2039), .D(n1807), 
        .Q(readOutBus[769]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_130_ ( .G(n2039), .D(n1809), 
        .Q(readOutBus[770]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_131_ ( .G(n2039), .D(n1811), 
        .Q(readOutBus[771]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_136_ ( .G(n2037), .D(n1821), 
        .Q(readOutBus[776]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_137_ ( .G(n2037), .D(n1823), 
        .Q(readOutBus[777]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_138_ ( .G(n2037), .D(n1825), 
        .Q(readOutBus[778]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_139_ ( .G(n2037), .D(n1827), 
        .Q(readOutBus[779]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_140_ ( .G(n2036), .D(n1829), 
        .Q(readOutBus[780]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_141_ ( .G(n2036), .D(n1831), 
        .Q(readOutBus[781]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_142_ ( .G(n2036), .D(n1833), 
        .Q(readOutBus[782]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_143_ ( .G(n2036), .D(n1835), 
        .Q(readOutBus[783]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_156_ ( .G(n2032), .D(n1861), 
        .Q(readOutBus[796]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_157_ ( .G(n2032), .D(n1863), 
        .Q(readOutBus[797]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_158_ ( .G(n2032), .D(n1865), 
        .Q(readOutBus[798]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_159_ ( .G(n2032), .D(n1867), 
        .Q(readOutBus[799]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_0_ ( .G(n1917), .D(n1549), 
        .Q(readOutBus[0]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_1_ ( .G(n1917), .D(n1551), 
        .Q(readOutBus[1]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_2_ ( .G(n1917), .D(n1553), 
        .Q(readOutBus[2]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_3_ ( .G(n1917), .D(n1555), 
        .Q(readOutBus[3]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_8_ ( .G(n1916), .D(n1565), 
        .Q(readOutBus[8]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_9_ ( .G(n1916), .D(n1567), 
        .Q(readOutBus[9]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_10_ ( .G(n1916), .D(n1569), 
        .Q(readOutBus[10]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_11_ ( .G(n1916), .D(n1571), 
        .Q(readOutBus[11]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_36_ ( .G(n1909), .D(n1621), 
        .Q(readOutBus[36]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_37_ ( .G(n1909), .D(n1623), 
        .Q(readOutBus[37]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_38_ ( .G(n1909), .D(n1625), 
        .Q(readOutBus[38]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_39_ ( .G(n1909), .D(n1627), 
        .Q(readOutBus[39]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_80_ ( .G(n1898), .D(n1709), 
        .Q(readOutBus[80]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_81_ ( .G(n1898), .D(n1711), 
        .Q(readOutBus[81]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_82_ ( .G(n1898), .D(n1713), 
        .Q(readOutBus[82]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_83_ ( .G(n1898), .D(n1715), 
        .Q(readOutBus[83]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_108_ ( .G(n1891), .D(n1765), 
        .Q(readOutBus[108]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_109_ ( .G(n1891), .D(n1767), 
        .Q(readOutBus[109]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_110_ ( .G(n1891), .D(n1769), 
        .Q(readOutBus[110]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_111_ ( .G(n1891), .D(n1771), 
        .Q(readOutBus[111]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_116_ ( .G(n1889), .D(n1781), 
        .Q(readOutBus[116]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_117_ ( .G(n1889), .D(n1783), 
        .Q(readOutBus[117]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_118_ ( .G(n1889), .D(n1785), 
        .Q(readOutBus[118]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_119_ ( .G(n1889), .D(n1787), 
        .Q(readOutBus[119]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_148_ ( .G(n1882), .D(n1845), 
        .Q(readOutBus[148]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_149_ ( .G(n1882), .D(n1847), 
        .Q(readOutBus[149]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_150_ ( .G(n1882), .D(n1849), 
        .Q(readOutBus[150]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_151_ ( .G(n1882), .D(n1851), 
        .Q(readOutBus[151]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_0_ ( .G(n1993), .D(n1549), 
        .Q(readOutBus[320]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_1_ ( .G(n1993), .D(n1551), 
        .Q(readOutBus[321]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_2_ ( .G(n1993), .D(n1553), 
        .Q(readOutBus[322]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_3_ ( .G(n1993), .D(n1555), 
        .Q(readOutBus[323]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_8_ ( .G(n1992), .D(n1565), 
        .Q(readOutBus[328]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_9_ ( .G(n1992), .D(n1567), 
        .Q(readOutBus[329]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_10_ ( .G(n1992), .D(n1569), 
        .Q(readOutBus[330]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_11_ ( .G(n1992), .D(n1571), 
        .Q(readOutBus[331]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_36_ ( .G(n1985), .D(n1621), 
        .Q(readOutBus[356]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_37_ ( .G(n1985), .D(n1623), 
        .Q(readOutBus[357]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_38_ ( .G(n1985), .D(n1625), 
        .Q(readOutBus[358]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_39_ ( .G(n1985), .D(n1627), 
        .Q(readOutBus[359]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_80_ ( .G(n1974), .D(n1709), 
        .Q(readOutBus[400]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_81_ ( .G(n1974), .D(n1711), 
        .Q(readOutBus[401]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_82_ ( .G(n1974), .D(n1713), 
        .Q(readOutBus[402]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_83_ ( .G(n1974), .D(n1715), 
        .Q(readOutBus[403]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_108_ ( .G(n1967), .D(n1765), 
        .Q(readOutBus[428]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_109_ ( .G(n1967), .D(n1767), 
        .Q(readOutBus[429]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_110_ ( .G(n1967), .D(n1769), 
        .Q(readOutBus[430]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_111_ ( .G(n1967), .D(n1771), 
        .Q(readOutBus[431]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_116_ ( .G(n1965), .D(n1781), 
        .Q(readOutBus[436]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_117_ ( .G(n1965), .D(n1783), 
        .Q(readOutBus[437]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_118_ ( .G(n1965), .D(n1785), 
        .Q(readOutBus[438]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_119_ ( .G(n1965), .D(n1787), 
        .Q(readOutBus[439]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_148_ ( .G(n1958), .D(n1845), 
        .Q(readOutBus[468]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_149_ ( .G(n1958), .D(n1847), 
        .Q(readOutBus[469]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_150_ ( .G(n1958), .D(n1849), 
        .Q(readOutBus[470]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_151_ ( .G(n1958), .D(n1851), 
        .Q(readOutBus[471]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_0_ ( .G(n2069), .D(n1549), 
        .Q(readOutBus[640]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_1_ ( .G(n2069), .D(n1551), 
        .Q(readOutBus[641]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_2_ ( .G(n2069), .D(n1553), 
        .Q(readOutBus[642]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_3_ ( .G(n2069), .D(n1555), 
        .Q(readOutBus[643]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_8_ ( .G(n2068), .D(n1565), 
        .Q(readOutBus[648]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_9_ ( .G(n2068), .D(n1567), 
        .Q(readOutBus[649]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_10_ ( .G(n2068), .D(n1569), 
        .Q(readOutBus[650]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_11_ ( .G(n2068), .D(n1571), 
        .Q(readOutBus[651]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_36_ ( .G(n2061), .D(n1621), 
        .Q(readOutBus[676]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_37_ ( .G(n2061), .D(n1623), 
        .Q(readOutBus[677]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_38_ ( .G(n2061), .D(n1625), 
        .Q(readOutBus[678]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_39_ ( .G(n2061), .D(n1627), 
        .Q(readOutBus[679]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_80_ ( .G(n2050), .D(n1709), 
        .Q(readOutBus[720]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_81_ ( .G(n2050), .D(n1711), 
        .Q(readOutBus[721]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_82_ ( .G(n2050), .D(n1713), 
        .Q(readOutBus[722]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_83_ ( .G(n2050), .D(n1715), 
        .Q(readOutBus[723]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_108_ ( .G(n2043), .D(n1765), 
        .Q(readOutBus[748]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_109_ ( .G(n2043), .D(n1767), 
        .Q(readOutBus[749]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_110_ ( .G(n2043), .D(n1769), 
        .Q(readOutBus[750]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_111_ ( .G(n2043), .D(n1771), 
        .Q(readOutBus[751]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_116_ ( .G(n2041), .D(n1781), 
        .Q(readOutBus[756]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_117_ ( .G(n2041), .D(n1783), 
        .Q(readOutBus[757]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_118_ ( .G(n2041), .D(n1785), 
        .Q(readOutBus[758]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_119_ ( .G(n2041), .D(n1787), 
        .Q(readOutBus[759]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_148_ ( .G(n2034), .D(n1845), 
        .Q(readOutBus[788]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_149_ ( .G(n2034), .D(n1847), 
        .Q(readOutBus[789]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_150_ ( .G(n2034), .D(n1849), 
        .Q(readOutBus[790]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_151_ ( .G(n2034), .D(n1851), 
        .Q(readOutBus[791]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_152_ ( .G(n2033), .D(n1853), 
        .Q(readOutBus[792]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_153_ ( .G(n2033), .D(n1855), 
        .Q(readOutBus[793]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_154_ ( .G(n2033), .D(n1857), 
        .Q(readOutBus[794]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_155_ ( .G(n2033), .D(n1859), 
        .Q(readOutBus[795]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_12_ ( .G(n1915), .D(n1573), 
        .Q(readOutBus[12]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_13_ ( .G(n1915), .D(n1575), 
        .Q(readOutBus[13]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_14_ ( .G(n1915), .D(n1577), 
        .Q(readOutBus[14]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_15_ ( .G(n1915), .D(n1579), 
        .Q(readOutBus[15]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_16_ ( .G(n1914), .D(n1581), 
        .Q(readOutBus[16]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_17_ ( .G(n1914), .D(n1583), 
        .Q(readOutBus[17]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_18_ ( .G(n1914), .D(n1585), 
        .Q(readOutBus[18]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_19_ ( .G(n1914), .D(n1587), 
        .Q(readOutBus[19]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_20_ ( .G(n1913), .D(n1589), 
        .Q(readOutBus[20]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_21_ ( .G(n1913), .D(n1591), 
        .Q(readOutBus[21]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_22_ ( .G(n1913), .D(n1593), 
        .Q(readOutBus[22]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_23_ ( .G(n1913), .D(n1595), 
        .Q(readOutBus[23]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_24_ ( .G(n1912), .D(n1597), 
        .Q(readOutBus[24]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_25_ ( .G(n1912), .D(n1599), 
        .Q(readOutBus[25]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_26_ ( .G(n1912), .D(n1601), 
        .Q(readOutBus[26]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_27_ ( .G(n1912), .D(n1603), 
        .Q(readOutBus[27]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_28_ ( .G(n1911), .D(n1605), 
        .Q(readOutBus[28]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_29_ ( .G(n1911), .D(n1607), 
        .Q(readOutBus[29]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_30_ ( .G(n1911), .D(n1609), 
        .Q(readOutBus[30]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_31_ ( .G(n1911), .D(n1611), 
        .Q(readOutBus[31]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_32_ ( .G(n1910), .D(n1613), 
        .Q(readOutBus[32]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_33_ ( .G(n1910), .D(n1615), 
        .Q(readOutBus[33]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_34_ ( .G(n1910), .D(n1617), 
        .Q(readOutBus[34]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_35_ ( .G(n1910), .D(n1619), 
        .Q(readOutBus[35]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_40_ ( .G(n1908), .D(n1629), 
        .Q(readOutBus[40]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_41_ ( .G(n1908), .D(n1631), 
        .Q(readOutBus[41]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_42_ ( .G(n1908), .D(n1633), 
        .Q(readOutBus[42]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_43_ ( .G(n1908), .D(n1635), 
        .Q(readOutBus[43]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_48_ ( .G(n1906), .D(n1645), 
        .Q(readOutBus[48]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_49_ ( .G(n1906), .D(n1647), 
        .Q(readOutBus[49]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_50_ ( .G(n1906), .D(n1649), 
        .Q(readOutBus[50]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_51_ ( .G(n1906), .D(n1651), 
        .Q(readOutBus[51]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_52_ ( .G(n1905), .D(n1653), 
        .Q(readOutBus[52]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_53_ ( .G(n1905), .D(n1655), 
        .Q(readOutBus[53]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_54_ ( .G(n1905), .D(n1657), 
        .Q(readOutBus[54]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_55_ ( .G(n1905), .D(n1659), 
        .Q(readOutBus[55]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_56_ ( .G(n1904), .D(n1661), 
        .Q(readOutBus[56]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_57_ ( .G(n1904), .D(n1663), 
        .Q(readOutBus[57]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_58_ ( .G(n1904), .D(n1665), 
        .Q(readOutBus[58]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_59_ ( .G(n1904), .D(n1667), 
        .Q(readOutBus[59]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_60_ ( .G(n1903), .D(n1669), 
        .Q(readOutBus[60]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_61_ ( .G(n1903), .D(n1671), 
        .Q(readOutBus[61]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_62_ ( .G(n1903), .D(n1673), 
        .Q(readOutBus[62]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_63_ ( .G(n1903), .D(n1675), 
        .Q(readOutBus[63]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_64_ ( .G(n1902), .D(n1677), 
        .Q(readOutBus[64]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_65_ ( .G(n1902), .D(n1679), 
        .Q(readOutBus[65]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_66_ ( .G(n1902), .D(n1681), 
        .Q(readOutBus[66]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_67_ ( .G(n1902), .D(n1683), 
        .Q(readOutBus[67]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_68_ ( .G(n1901), .D(n1685), 
        .Q(readOutBus[68]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_69_ ( .G(n1901), .D(n1687), 
        .Q(readOutBus[69]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_70_ ( .G(n1901), .D(n1689), 
        .Q(readOutBus[70]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_71_ ( .G(n1901), .D(n1691), 
        .Q(readOutBus[71]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_72_ ( .G(n1900), .D(n1693), 
        .Q(readOutBus[72]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_73_ ( .G(n1900), .D(n1695), 
        .Q(readOutBus[73]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_74_ ( .G(n1900), .D(n1697), 
        .Q(readOutBus[74]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_75_ ( .G(n1900), .D(n1699), 
        .Q(readOutBus[75]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_96_ ( .G(n1894), .D(n1741), 
        .Q(readOutBus[96]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_97_ ( .G(n1894), .D(n1743), 
        .Q(readOutBus[97]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_98_ ( .G(n1894), .D(n1745), 
        .Q(readOutBus[98]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_99_ ( .G(n1894), .D(n1747), 
        .Q(readOutBus[99]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_100_ ( .G(n1893), .D(n1749), 
        .Q(readOutBus[100]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_101_ ( .G(n1893), .D(n1751), 
        .Q(readOutBus[101]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_102_ ( .G(n1893), .D(n1753), 
        .Q(readOutBus[102]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_103_ ( .G(n1893), .D(n1755), 
        .Q(readOutBus[103]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_104_ ( .G(n1892), .D(n1757), 
        .Q(readOutBus[104]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_105_ ( .G(n1892), .D(n1759), 
        .Q(readOutBus[105]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_106_ ( .G(n1892), .D(n1761), 
        .Q(readOutBus[106]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_107_ ( .G(n1892), .D(n1763), 
        .Q(readOutBus[107]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_112_ ( .G(n1890), .D(n1773), 
        .Q(readOutBus[112]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_113_ ( .G(n1890), .D(n1775), 
        .Q(readOutBus[113]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_114_ ( .G(n1890), .D(n1777), 
        .Q(readOutBus[114]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_115_ ( .G(n1890), .D(n1779), 
        .Q(readOutBus[115]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_12_ ( .G(n1991), .D(n1573), 
        .Q(readOutBus[332]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_13_ ( .G(n1991), .D(n1575), 
        .Q(readOutBus[333]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_14_ ( .G(n1991), .D(n1577), 
        .Q(readOutBus[334]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_15_ ( .G(n1991), .D(n1579), 
        .Q(readOutBus[335]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_16_ ( .G(n1990), .D(n1581), 
        .Q(readOutBus[336]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_17_ ( .G(n1990), .D(n1583), 
        .Q(readOutBus[337]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_18_ ( .G(n1990), .D(n1585), 
        .Q(readOutBus[338]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_19_ ( .G(n1990), .D(n1587), 
        .Q(readOutBus[339]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_20_ ( .G(n1989), .D(n1589), 
        .Q(readOutBus[340]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_21_ ( .G(n1989), .D(n1591), 
        .Q(readOutBus[341]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_22_ ( .G(n1989), .D(n1593), 
        .Q(readOutBus[342]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_23_ ( .G(n1989), .D(n1595), 
        .Q(readOutBus[343]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_24_ ( .G(n1988), .D(n1597), 
        .Q(readOutBus[344]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_25_ ( .G(n1988), .D(n1599), 
        .Q(readOutBus[345]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_26_ ( .G(n1988), .D(n1601), 
        .Q(readOutBus[346]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_27_ ( .G(n1988), .D(n1603), 
        .Q(readOutBus[347]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_28_ ( .G(n1987), .D(n1605), 
        .Q(readOutBus[348]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_29_ ( .G(n1987), .D(n1607), 
        .Q(readOutBus[349]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_30_ ( .G(n1987), .D(n1609), 
        .Q(readOutBus[350]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_31_ ( .G(n1987), .D(n1611), 
        .Q(readOutBus[351]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_32_ ( .G(n1986), .D(n1613), 
        .Q(readOutBus[352]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_33_ ( .G(n1986), .D(n1615), 
        .Q(readOutBus[353]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_34_ ( .G(n1986), .D(n1617), 
        .Q(readOutBus[354]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_35_ ( .G(n1986), .D(n1619), 
        .Q(readOutBus[355]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_40_ ( .G(n1984), .D(n1629), 
        .Q(readOutBus[360]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_41_ ( .G(n1984), .D(n1631), 
        .Q(readOutBus[361]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_42_ ( .G(n1984), .D(n1633), 
        .Q(readOutBus[362]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_43_ ( .G(n1984), .D(n1635), 
        .Q(readOutBus[363]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_48_ ( .G(n1982), .D(n1645), 
        .Q(readOutBus[368]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_49_ ( .G(n1982), .D(n1647), 
        .Q(readOutBus[369]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_50_ ( .G(n1982), .D(n1649), 
        .Q(readOutBus[370]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_51_ ( .G(n1982), .D(n1651), 
        .Q(readOutBus[371]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_52_ ( .G(n1981), .D(n1653), 
        .Q(readOutBus[372]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_53_ ( .G(n1981), .D(n1655), 
        .Q(readOutBus[373]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_54_ ( .G(n1981), .D(n1657), 
        .Q(readOutBus[374]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_55_ ( .G(n1981), .D(n1659), 
        .Q(readOutBus[375]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_56_ ( .G(n1980), .D(n1661), 
        .Q(readOutBus[376]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_57_ ( .G(n1980), .D(n1663), 
        .Q(readOutBus[377]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_58_ ( .G(n1980), .D(n1665), 
        .Q(readOutBus[378]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_59_ ( .G(n1980), .D(n1667), 
        .Q(readOutBus[379]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_60_ ( .G(n1979), .D(n1669), 
        .Q(readOutBus[380]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_61_ ( .G(n1979), .D(n1671), 
        .Q(readOutBus[381]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_62_ ( .G(n1979), .D(n1673), 
        .Q(readOutBus[382]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_63_ ( .G(n1979), .D(n1675), 
        .Q(readOutBus[383]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_64_ ( .G(n1978), .D(n1677), 
        .Q(readOutBus[384]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_65_ ( .G(n1978), .D(n1679), 
        .Q(readOutBus[385]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_66_ ( .G(n1978), .D(n1681), 
        .Q(readOutBus[386]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_67_ ( .G(n1978), .D(n1683), 
        .Q(readOutBus[387]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_68_ ( .G(n1977), .D(n1685), 
        .Q(readOutBus[388]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_69_ ( .G(n1977), .D(n1687), 
        .Q(readOutBus[389]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_70_ ( .G(n1977), .D(n1689), 
        .Q(readOutBus[390]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_71_ ( .G(n1977), .D(n1691), 
        .Q(readOutBus[391]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_72_ ( .G(n1976), .D(n1693), 
        .Q(readOutBus[392]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_73_ ( .G(n1976), .D(n1695), 
        .Q(readOutBus[393]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_74_ ( .G(n1976), .D(n1697), 
        .Q(readOutBus[394]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_75_ ( .G(n1976), .D(n1699), 
        .Q(readOutBus[395]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_96_ ( .G(n1970), .D(n1741), 
        .Q(readOutBus[416]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_97_ ( .G(n1970), .D(n1743), 
        .Q(readOutBus[417]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_98_ ( .G(n1970), .D(n1745), 
        .Q(readOutBus[418]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_99_ ( .G(n1970), .D(n1747), 
        .Q(readOutBus[419]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_100_ ( .G(n1969), .D(n1749), 
        .Q(readOutBus[420]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_101_ ( .G(n1969), .D(n1751), 
        .Q(readOutBus[421]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_102_ ( .G(n1969), .D(n1753), 
        .Q(readOutBus[422]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_103_ ( .G(n1969), .D(n1755), 
        .Q(readOutBus[423]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_104_ ( .G(n1968), .D(n1757), 
        .Q(readOutBus[424]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_105_ ( .G(n1968), .D(n1759), 
        .Q(readOutBus[425]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_106_ ( .G(n1968), .D(n1761), 
        .Q(readOutBus[426]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_107_ ( .G(n1968), .D(n1763), 
        .Q(readOutBus[427]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_112_ ( .G(n1966), .D(n1773), 
        .Q(readOutBus[432]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_113_ ( .G(n1966), .D(n1775), 
        .Q(readOutBus[433]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_114_ ( .G(n1966), .D(n1777), 
        .Q(readOutBus[434]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_115_ ( .G(n1966), .D(n1779), 
        .Q(readOutBus[435]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_12_ ( .G(n2067), .D(n1573), 
        .Q(readOutBus[652]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_13_ ( .G(n2067), .D(n1575), 
        .Q(readOutBus[653]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_14_ ( .G(n2067), .D(n1577), 
        .Q(readOutBus[654]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_15_ ( .G(n2067), .D(n1579), 
        .Q(readOutBus[655]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_16_ ( .G(n2066), .D(n1581), 
        .Q(readOutBus[656]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_17_ ( .G(n2066), .D(n1583), 
        .Q(readOutBus[657]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_18_ ( .G(n2066), .D(n1585), 
        .Q(readOutBus[658]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_19_ ( .G(n2066), .D(n1587), 
        .Q(readOutBus[659]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_20_ ( .G(n2065), .D(n1589), 
        .Q(readOutBus[660]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_21_ ( .G(n2065), .D(n1591), 
        .Q(readOutBus[661]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_22_ ( .G(n2065), .D(n1593), 
        .Q(readOutBus[662]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_23_ ( .G(n2065), .D(n1595), 
        .Q(readOutBus[663]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_24_ ( .G(n2064), .D(n1597), 
        .Q(readOutBus[664]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_25_ ( .G(n2064), .D(n1599), 
        .Q(readOutBus[665]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_26_ ( .G(n2064), .D(n1601), 
        .Q(readOutBus[666]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_27_ ( .G(n2064), .D(n1603), 
        .Q(readOutBus[667]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_28_ ( .G(n2063), .D(n1605), 
        .Q(readOutBus[668]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_29_ ( .G(n2063), .D(n1607), 
        .Q(readOutBus[669]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_30_ ( .G(n2063), .D(n1609), 
        .Q(readOutBus[670]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_31_ ( .G(n2063), .D(n1611), 
        .Q(readOutBus[671]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_32_ ( .G(n2062), .D(n1613), 
        .Q(readOutBus[672]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_33_ ( .G(n2062), .D(n1615), 
        .Q(readOutBus[673]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_34_ ( .G(n2062), .D(n1617), 
        .Q(readOutBus[674]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_35_ ( .G(n2062), .D(n1619), 
        .Q(readOutBus[675]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_40_ ( .G(n2060), .D(n1629), 
        .Q(readOutBus[680]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_41_ ( .G(n2060), .D(n1631), 
        .Q(readOutBus[681]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_42_ ( .G(n2060), .D(n1633), 
        .Q(readOutBus[682]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_43_ ( .G(n2060), .D(n1635), 
        .Q(readOutBus[683]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_48_ ( .G(n2058), .D(n1645), 
        .Q(readOutBus[688]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_49_ ( .G(n2058), .D(n1647), 
        .Q(readOutBus[689]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_50_ ( .G(n2058), .D(n1649), 
        .Q(readOutBus[690]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_51_ ( .G(n2058), .D(n1651), 
        .Q(readOutBus[691]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_52_ ( .G(n2057), .D(n1653), 
        .Q(readOutBus[692]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_53_ ( .G(n2057), .D(n1655), 
        .Q(readOutBus[693]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_54_ ( .G(n2057), .D(n1657), 
        .Q(readOutBus[694]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_55_ ( .G(n2057), .D(n1659), 
        .Q(readOutBus[695]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_56_ ( .G(n2056), .D(n1661), 
        .Q(readOutBus[696]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_57_ ( .G(n2056), .D(n1663), 
        .Q(readOutBus[697]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_58_ ( .G(n2056), .D(n1665), 
        .Q(readOutBus[698]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_59_ ( .G(n2056), .D(n1667), 
        .Q(readOutBus[699]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_60_ ( .G(n2055), .D(n1669), 
        .Q(readOutBus[700]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_61_ ( .G(n2055), .D(n1671), 
        .Q(readOutBus[701]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_62_ ( .G(n2055), .D(n1673), 
        .Q(readOutBus[702]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_63_ ( .G(n2055), .D(n1675), 
        .Q(readOutBus[703]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_64_ ( .G(n2054), .D(n1677), 
        .Q(readOutBus[704]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_65_ ( .G(n2054), .D(n1679), 
        .Q(readOutBus[705]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_66_ ( .G(n2054), .D(n1681), 
        .Q(readOutBus[706]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_67_ ( .G(n2054), .D(n1683), 
        .Q(readOutBus[707]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_68_ ( .G(n2053), .D(n1685), 
        .Q(readOutBus[708]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_69_ ( .G(n2053), .D(n1687), 
        .Q(readOutBus[709]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_70_ ( .G(n2053), .D(n1689), 
        .Q(readOutBus[710]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_71_ ( .G(n2053), .D(n1691), 
        .Q(readOutBus[711]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_72_ ( .G(n2052), .D(n1693), 
        .Q(readOutBus[712]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_73_ ( .G(n2052), .D(n1695), 
        .Q(readOutBus[713]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_74_ ( .G(n2052), .D(n1697), 
        .Q(readOutBus[714]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_75_ ( .G(n2052), .D(n1699), 
        .Q(readOutBus[715]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_96_ ( .G(n2046), .D(n1741), 
        .Q(readOutBus[736]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_97_ ( .G(n2046), .D(n1743), 
        .Q(readOutBus[737]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_98_ ( .G(n2046), .D(n1745), 
        .Q(readOutBus[738]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_99_ ( .G(n2046), .D(n1747), 
        .Q(readOutBus[739]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_100_ ( .G(n2045), .D(n1749), 
        .Q(readOutBus[740]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_101_ ( .G(n2045), .D(n1751), 
        .Q(readOutBus[741]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_102_ ( .G(n2045), .D(n1753), 
        .Q(readOutBus[742]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_103_ ( .G(n2045), .D(n1755), 
        .Q(readOutBus[743]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_104_ ( .G(n2044), .D(n1757), 
        .Q(readOutBus[744]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_105_ ( .G(n2044), .D(n1759), 
        .Q(readOutBus[745]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_106_ ( .G(n2044), .D(n1761), 
        .Q(readOutBus[746]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_107_ ( .G(n2044), .D(n1763), 
        .Q(readOutBus[747]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_112_ ( .G(n2042), .D(n1773), 
        .Q(readOutBus[752]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_113_ ( .G(n2042), .D(n1775), 
        .Q(readOutBus[753]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_114_ ( .G(n2042), .D(n1777), 
        .Q(readOutBus[754]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_115_ ( .G(n2042), .D(n1779), 
        .Q(readOutBus[755]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_144_ ( .G(n2035), .D(n1837), 
        .Q(readOutBus[784]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_145_ ( .G(n2035), .D(n1839), 
        .Q(readOutBus[785]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_146_ ( .G(n2035), .D(n1841), 
        .Q(readOutBus[786]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_147_ ( .G(n2035), .D(n1843), 
        .Q(readOutBus[787]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_132_ ( .G(n2038), .D(n1813), 
        .Q(readOutBus[772]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_133_ ( .G(n2038), .D(n1815), 
        .Q(readOutBus[773]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_134_ ( .G(n2038), .D(n1817), 
        .Q(readOutBus[774]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_135_ ( .G(n2038), .D(n1819), 
        .Q(readOutBus[775]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_5_ ( .G(n1868), .D(n1559), 
        .Q(readOutBus[5]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_7_ ( .G(n1868), .D(n1563), 
        .Q(readOutBus[7]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_5_ ( .G(n1872), .D(n1559), 
        .Q(readOutBus[325]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_7_ ( .G(n1872), .D(n1563), 
        .Q(readOutBus[327]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_5_ ( .G(n1876), .D(n1559), 
        .Q(readOutBus[645]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_7_ ( .G(n1876), .D(n1563), 
        .Q(readOutBus[647]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_4_ ( .G(n1869), .D(n1557), 
        .Q(readOutBus[4]) );
  TLATXLTS Generate_Node_Banks_0__NB_readOut_reg_6_ ( .G(n1869), .D(n1561), 
        .Q(readOutBus[6]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_4_ ( .G(n1873), .D(n1557), 
        .Q(readOutBus[324]) );
  TLATXLTS Generate_Node_Banks_2__NB_readOut_reg_6_ ( .G(n1873), .D(n1561), 
        .Q(readOutBus[326]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_4_ ( .G(n1877), .D(n1557), 
        .Q(readOutBus[644]) );
  TLATXLTS Generate_Node_Banks_4__NB_readOut_reg_6_ ( .G(n1877), .D(n1561), 
        .Q(readOutBus[646]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_44_ ( .G(n1945), .D(n1636), 
        .Q(readOutBus[204]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_45_ ( .G(n1945), .D(n1638), 
        .Q(readOutBus[205]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_46_ ( .G(n1945), .D(n1640), 
        .Q(readOutBus[206]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_47_ ( .G(n1945), .D(n1642), 
        .Q(readOutBus[207]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_76_ ( .G(n1937), .D(n1700), 
        .Q(readOutBus[236]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_77_ ( .G(n1937), .D(n1702), 
        .Q(readOutBus[237]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_78_ ( .G(n1937), .D(n1704), 
        .Q(readOutBus[238]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_79_ ( .G(n1937), .D(n1706), 
        .Q(readOutBus[239]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_84_ ( .G(n1935), .D(n1716), 
        .Q(readOutBus[244]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_85_ ( .G(n1935), .D(n1718), 
        .Q(readOutBus[245]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_86_ ( .G(n1935), .D(n1720), 
        .Q(readOutBus[246]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_87_ ( .G(n1935), .D(n1722), 
        .Q(readOutBus[247]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_88_ ( .G(n1934), .D(n1724), 
        .Q(readOutBus[248]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_89_ ( .G(n1934), .D(n1726), 
        .Q(readOutBus[249]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_90_ ( .G(n1934), .D(n1728), 
        .Q(readOutBus[250]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_91_ ( .G(n1934), .D(n1730), 
        .Q(readOutBus[251]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_92_ ( .G(n1933), .D(n1732), 
        .Q(readOutBus[252]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_93_ ( .G(n1933), .D(n1734), 
        .Q(readOutBus[253]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_94_ ( .G(n1933), .D(n1736), 
        .Q(readOutBus[254]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_95_ ( .G(n1933), .D(n1738), 
        .Q(readOutBus[255]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_120_ ( .G(n738), .D(n1788), 
        .Q(readOutBus[280]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_121_ ( .G(n739), .D(n1790), 
        .Q(readOutBus[281]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_122_ ( .G(n717), .D(n1792), 
        .Q(readOutBus[282]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_123_ ( .G(n719), .D(n1794), 
        .Q(readOutBus[283]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_124_ ( .G(n1926), .D(n1796), 
        .Q(readOutBus[284]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_125_ ( .G(n1926), .D(n1798), 
        .Q(readOutBus[285]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_126_ ( .G(n1926), .D(n1800), 
        .Q(readOutBus[286]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_127_ ( .G(n1926), .D(n1802), 
        .Q(readOutBus[287]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_128_ ( .G(n1925), .D(n1804), 
        .Q(readOutBus[288]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_129_ ( .G(n1925), .D(n1806), 
        .Q(readOutBus[289]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_130_ ( .G(n1925), .D(n1808), 
        .Q(readOutBus[290]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_131_ ( .G(n1925), .D(n1810), 
        .Q(readOutBus[291]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_132_ ( .G(n1924), .D(n1812), 
        .Q(readOutBus[292]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_133_ ( .G(n1924), .D(n1814), 
        .Q(readOutBus[293]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_134_ ( .G(n1924), .D(n1816), 
        .Q(readOutBus[294]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_135_ ( .G(n1924), .D(n1818), 
        .Q(readOutBus[295]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_136_ ( .G(n1923), .D(n1820), 
        .Q(readOutBus[296]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_137_ ( .G(n1923), .D(n1822), 
        .Q(readOutBus[297]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_138_ ( .G(n1923), .D(n1824), 
        .Q(readOutBus[298]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_139_ ( .G(n1923), .D(n1826), 
        .Q(readOutBus[299]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_140_ ( .G(n1922), .D(n1828), 
        .Q(readOutBus[300]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_141_ ( .G(n1922), .D(n1830), 
        .Q(readOutBus[301]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_142_ ( .G(n1922), .D(n1832), 
        .Q(readOutBus[302]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_143_ ( .G(n1922), .D(n1834), 
        .Q(readOutBus[303]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_144_ ( .G(n1921), .D(n1836), 
        .Q(readOutBus[304]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_145_ ( .G(n1921), .D(n1838), 
        .Q(readOutBus[305]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_146_ ( .G(n1921), .D(n1840), 
        .Q(readOutBus[306]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_147_ ( .G(n1921), .D(n1842), 
        .Q(readOutBus[307]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_152_ ( .G(n1919), .D(n1852), 
        .Q(readOutBus[312]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_153_ ( .G(n1919), .D(n1854), 
        .Q(readOutBus[313]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_154_ ( .G(n1919), .D(n1856), 
        .Q(readOutBus[314]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_155_ ( .G(n1919), .D(n1858), 
        .Q(readOutBus[315]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_156_ ( .G(n1918), .D(n1860), 
        .Q(readOutBus[316]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_44_ ( .G(n2021), .D(n1636), 
        .Q(readOutBus[524]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_45_ ( .G(n2021), .D(n1638), 
        .Q(readOutBus[525]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_46_ ( .G(n2021), .D(n1640), 
        .Q(readOutBus[526]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_47_ ( .G(n2021), .D(n1642), 
        .Q(readOutBus[527]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_76_ ( .G(n2013), .D(n1700), 
        .Q(readOutBus[556]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_77_ ( .G(n2013), .D(n1702), 
        .Q(readOutBus[557]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_78_ ( .G(n2013), .D(n1704), 
        .Q(readOutBus[558]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_79_ ( .G(n2013), .D(n1706), 
        .Q(readOutBus[559]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_84_ ( .G(n2011), .D(n1716), 
        .Q(readOutBus[564]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_85_ ( .G(n2011), .D(n1718), 
        .Q(readOutBus[565]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_86_ ( .G(n2011), .D(n1720), 
        .Q(readOutBus[566]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_87_ ( .G(n2011), .D(n1722), 
        .Q(readOutBus[567]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_88_ ( .G(n2010), .D(n1724), 
        .Q(readOutBus[568]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_89_ ( .G(n2010), .D(n1726), 
        .Q(readOutBus[569]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_90_ ( .G(n2010), .D(n1728), 
        .Q(readOutBus[570]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_91_ ( .G(n2010), .D(n1730), 
        .Q(readOutBus[571]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_92_ ( .G(n2009), .D(n1732), 
        .Q(readOutBus[572]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_93_ ( .G(n2009), .D(n1734), 
        .Q(readOutBus[573]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_94_ ( .G(n2009), .D(n1736), 
        .Q(readOutBus[574]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_95_ ( .G(n2009), .D(n1738), 
        .Q(readOutBus[575]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_120_ ( .G(n735), .D(n1788), 
        .Q(readOutBus[600]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_121_ ( .G(n736), .D(n1790), 
        .Q(readOutBus[601]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_122_ ( .G(n716), .D(n1792), 
        .Q(readOutBus[602]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_123_ ( .G(n718), .D(n1794), 
        .Q(readOutBus[603]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_124_ ( .G(n2002), .D(n1796), 
        .Q(readOutBus[604]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_125_ ( .G(n2002), .D(n1798), 
        .Q(readOutBus[605]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_126_ ( .G(n2002), .D(n1800), 
        .Q(readOutBus[606]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_127_ ( .G(n2002), .D(n1802), 
        .Q(readOutBus[607]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_128_ ( .G(n2001), .D(n1804), 
        .Q(readOutBus[608]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_129_ ( .G(n2001), .D(n1806), 
        .Q(readOutBus[609]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_130_ ( .G(n2001), .D(n1808), 
        .Q(readOutBus[610]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_131_ ( .G(n2001), .D(n1810), 
        .Q(readOutBus[611]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_132_ ( .G(n2000), .D(n1812), 
        .Q(readOutBus[612]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_133_ ( .G(n2000), .D(n1814), 
        .Q(readOutBus[613]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_134_ ( .G(n2000), .D(n1816), 
        .Q(readOutBus[614]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_135_ ( .G(n2000), .D(n1818), 
        .Q(readOutBus[615]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_136_ ( .G(n1999), .D(n1820), 
        .Q(readOutBus[616]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_137_ ( .G(n1999), .D(n1822), 
        .Q(readOutBus[617]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_138_ ( .G(n1999), .D(n1824), 
        .Q(readOutBus[618]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_139_ ( .G(n1999), .D(n1826), 
        .Q(readOutBus[619]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_140_ ( .G(n1998), .D(n1828), 
        .Q(readOutBus[620]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_141_ ( .G(n1998), .D(n1830), 
        .Q(readOutBus[621]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_142_ ( .G(n1998), .D(n1832), 
        .Q(readOutBus[622]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_143_ ( .G(n1998), .D(n1834), 
        .Q(readOutBus[623]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_144_ ( .G(n1997), .D(n1836), 
        .Q(readOutBus[624]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_145_ ( .G(n1997), .D(n1838), 
        .Q(readOutBus[625]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_146_ ( .G(n1997), .D(n1840), 
        .Q(readOutBus[626]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_147_ ( .G(n1997), .D(n1842), 
        .Q(readOutBus[627]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_152_ ( .G(n1995), .D(n1852), 
        .Q(readOutBus[632]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_153_ ( .G(n1995), .D(n1854), 
        .Q(readOutBus[633]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_154_ ( .G(n1995), .D(n1856), 
        .Q(readOutBus[634]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_155_ ( .G(n1995), .D(n1858), 
        .Q(readOutBus[635]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_44_ ( .G(n2097), .D(n1636), 
        .Q(readOutBus[844]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_45_ ( .G(n2097), .D(n1638), 
        .Q(readOutBus[845]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_46_ ( .G(n2097), .D(n1640), 
        .Q(readOutBus[846]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_47_ ( .G(n2097), .D(n1642), 
        .Q(readOutBus[847]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_76_ ( .G(n2089), .D(n1700), 
        .Q(readOutBus[876]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_77_ ( .G(n2089), .D(n1702), 
        .Q(readOutBus[877]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_78_ ( .G(n2089), .D(n1704), 
        .Q(readOutBus[878]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_79_ ( .G(n2089), .D(n1706), 
        .Q(readOutBus[879]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_84_ ( .G(n2087), .D(n1716), 
        .Q(readOutBus[884]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_85_ ( .G(n2087), .D(n1718), 
        .Q(readOutBus[885]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_86_ ( .G(n2087), .D(n1720), 
        .Q(readOutBus[886]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_87_ ( .G(n2087), .D(n1722), 
        .Q(readOutBus[887]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_88_ ( .G(n2086), .D(n1724), 
        .Q(readOutBus[888]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_89_ ( .G(n2086), .D(n1726), 
        .Q(readOutBus[889]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_90_ ( .G(n2086), .D(n1728), 
        .Q(readOutBus[890]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_91_ ( .G(n2086), .D(n1730), 
        .Q(readOutBus[891]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_92_ ( .G(n2085), .D(n1732), 
        .Q(readOutBus[892]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_93_ ( .G(n2085), .D(n1734), 
        .Q(readOutBus[893]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_94_ ( .G(n2085), .D(n1736), 
        .Q(readOutBus[894]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_95_ ( .G(n2085), .D(n1738), 
        .Q(readOutBus[895]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_120_ ( .G(n2078), .D(n1788), 
        .Q(readOutBus[920]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_121_ ( .G(n2078), .D(n1790), 
        .Q(readOutBus[921]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_122_ ( .G(n2078), .D(n1792), 
        .Q(readOutBus[922]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_123_ ( .G(n2078), .D(n1794), 
        .Q(readOutBus[923]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_124_ ( .G(n2077), .D(n1796), 
        .Q(readOutBus[924]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_125_ ( .G(n2077), .D(n1798), 
        .Q(readOutBus[925]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_126_ ( .G(n2077), .D(n1800), 
        .Q(readOutBus[926]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_127_ ( .G(n2077), .D(n1802), 
        .Q(readOutBus[927]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_128_ ( .G(n734), .D(n1804), 
        .Q(readOutBus[928]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_129_ ( .G(n701), .D(n1806), 
        .Q(readOutBus[929]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_130_ ( .G(n712), .D(n1808), 
        .Q(readOutBus[930]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_131_ ( .G(n713), .D(n1810), 
        .Q(readOutBus[931]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_24_ ( .G(n1950), .D(n1596), 
        .Q(readOutBus[184]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_25_ ( .G(n1950), .D(n1598), 
        .Q(readOutBus[185]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_26_ ( .G(n1950), .D(n1600), 
        .Q(readOutBus[186]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_27_ ( .G(n1950), .D(n1602), 
        .Q(readOutBus[187]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_28_ ( .G(n1949), .D(n1604), 
        .Q(readOutBus[188]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_29_ ( .G(n1949), .D(n1606), 
        .Q(readOutBus[189]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_30_ ( .G(n1949), .D(n1608), 
        .Q(readOutBus[190]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_31_ ( .G(n1949), .D(n1610), 
        .Q(readOutBus[191]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_32_ ( .G(n1948), .D(n1612), 
        .Q(readOutBus[192]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_33_ ( .G(n1948), .D(n1614), 
        .Q(readOutBus[193]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_34_ ( .G(n1948), .D(n1616), 
        .Q(readOutBus[194]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_35_ ( .G(n1948), .D(n1618), 
        .Q(readOutBus[195]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_40_ ( .G(n1946), .D(n1628), 
        .Q(readOutBus[200]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_41_ ( .G(n1946), .D(n1630), 
        .Q(readOutBus[201]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_42_ ( .G(n1946), .D(n1632), 
        .Q(readOutBus[202]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_43_ ( .G(n1946), .D(n1634), 
        .Q(readOutBus[203]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_60_ ( .G(n1941), .D(n1668), 
        .Q(readOutBus[220]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_61_ ( .G(n1941), .D(n1670), 
        .Q(readOutBus[221]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_62_ ( .G(n1941), .D(n1672), 
        .Q(readOutBus[222]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_63_ ( .G(n1941), .D(n1674), 
        .Q(readOutBus[223]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_64_ ( .G(n1940), .D(n1676), 
        .Q(readOutBus[224]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_65_ ( .G(n1940), .D(n1678), 
        .Q(readOutBus[225]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_66_ ( .G(n1940), .D(n1680), 
        .Q(readOutBus[226]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_67_ ( .G(n1940), .D(n1682), 
        .Q(readOutBus[227]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_68_ ( .G(n1939), .D(n1684), 
        .Q(readOutBus[228]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_69_ ( .G(n1939), .D(n1686), 
        .Q(readOutBus[229]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_70_ ( .G(n1939), .D(n1688), 
        .Q(readOutBus[230]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_71_ ( .G(n1939), .D(n1690), 
        .Q(readOutBus[231]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_72_ ( .G(n1938), .D(n1692), 
        .Q(readOutBus[232]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_73_ ( .G(n1938), .D(n1694), 
        .Q(readOutBus[233]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_74_ ( .G(n1938), .D(n1696), 
        .Q(readOutBus[234]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_75_ ( .G(n1938), .D(n1698), 
        .Q(readOutBus[235]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_96_ ( .G(n1932), .D(n1740), 
        .Q(readOutBus[256]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_97_ ( .G(n1932), .D(n1742), 
        .Q(readOutBus[257]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_98_ ( .G(n1932), .D(n1744), 
        .Q(readOutBus[258]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_99_ ( .G(n1932), .D(n1746), 
        .Q(readOutBus[259]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_100_ ( .G(n1931), .D(n1748), 
        .Q(readOutBus[260]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_101_ ( .G(n1931), .D(n1750), 
        .Q(readOutBus[261]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_102_ ( .G(n1931), .D(n1752), 
        .Q(readOutBus[262]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_103_ ( .G(n1931), .D(n1754), 
        .Q(readOutBus[263]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_104_ ( .G(n1930), .D(n1756), 
        .Q(readOutBus[264]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_105_ ( .G(n1930), .D(n1758), 
        .Q(readOutBus[265]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_106_ ( .G(n1930), .D(n1760), 
        .Q(readOutBus[266]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_107_ ( .G(n1930), .D(n1762), 
        .Q(readOutBus[267]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_112_ ( .G(n1928), .D(n1772), 
        .Q(readOutBus[272]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_113_ ( .G(n1928), .D(n1774), 
        .Q(readOutBus[273]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_114_ ( .G(n1928), .D(n1776), 
        .Q(readOutBus[274]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_115_ ( .G(n1928), .D(n1778), 
        .Q(readOutBus[275]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_157_ ( .G(n1918), .D(n1862), 
        .Q(readOutBus[317]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_158_ ( .G(n1918), .D(n1864), 
        .Q(readOutBus[318]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_159_ ( .G(n1918), .D(n1866), 
        .Q(readOutBus[319]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_24_ ( .G(n2026), .D(n1596), 
        .Q(readOutBus[504]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_25_ ( .G(n2026), .D(n1598), 
        .Q(readOutBus[505]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_26_ ( .G(n2026), .D(n1600), 
        .Q(readOutBus[506]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_27_ ( .G(n2026), .D(n1602), 
        .Q(readOutBus[507]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_28_ ( .G(n2025), .D(n1604), 
        .Q(readOutBus[508]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_29_ ( .G(n2025), .D(n1606), 
        .Q(readOutBus[509]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_30_ ( .G(n2025), .D(n1608), 
        .Q(readOutBus[510]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_31_ ( .G(n2025), .D(n1610), 
        .Q(readOutBus[511]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_32_ ( .G(n2024), .D(n1612), 
        .Q(readOutBus[512]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_33_ ( .G(n2024), .D(n1614), 
        .Q(readOutBus[513]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_34_ ( .G(n2024), .D(n1616), 
        .Q(readOutBus[514]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_35_ ( .G(n2024), .D(n1618), 
        .Q(readOutBus[515]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_40_ ( .G(n2022), .D(n1628), 
        .Q(readOutBus[520]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_41_ ( .G(n2022), .D(n1630), 
        .Q(readOutBus[521]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_42_ ( .G(n2022), .D(n1632), 
        .Q(readOutBus[522]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_43_ ( .G(n2022), .D(n1634), 
        .Q(readOutBus[523]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_60_ ( .G(n2017), .D(n1668), 
        .Q(readOutBus[540]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_61_ ( .G(n2017), .D(n1670), 
        .Q(readOutBus[541]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_62_ ( .G(n2017), .D(n1672), 
        .Q(readOutBus[542]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_63_ ( .G(n2017), .D(n1674), 
        .Q(readOutBus[543]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_64_ ( .G(n2016), .D(n1676), 
        .Q(readOutBus[544]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_65_ ( .G(n2016), .D(n1678), 
        .Q(readOutBus[545]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_66_ ( .G(n2016), .D(n1680), 
        .Q(readOutBus[546]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_67_ ( .G(n2016), .D(n1682), 
        .Q(readOutBus[547]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_68_ ( .G(n2015), .D(n1684), 
        .Q(readOutBus[548]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_69_ ( .G(n2015), .D(n1686), 
        .Q(readOutBus[549]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_70_ ( .G(n2015), .D(n1688), 
        .Q(readOutBus[550]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_71_ ( .G(n2015), .D(n1690), 
        .Q(readOutBus[551]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_72_ ( .G(n2014), .D(n1692), 
        .Q(readOutBus[552]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_73_ ( .G(n2014), .D(n1694), 
        .Q(readOutBus[553]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_74_ ( .G(n2014), .D(n1696), 
        .Q(readOutBus[554]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_75_ ( .G(n2014), .D(n1698), 
        .Q(readOutBus[555]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_96_ ( .G(n2008), .D(n1740), 
        .Q(readOutBus[576]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_97_ ( .G(n2008), .D(n1742), 
        .Q(readOutBus[577]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_98_ ( .G(n2008), .D(n1744), 
        .Q(readOutBus[578]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_99_ ( .G(n2008), .D(n1746), 
        .Q(readOutBus[579]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_100_ ( .G(n2007), .D(n1748), 
        .Q(readOutBus[580]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_101_ ( .G(n2007), .D(n1750), 
        .Q(readOutBus[581]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_102_ ( .G(n2007), .D(n1752), 
        .Q(readOutBus[582]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_103_ ( .G(n2007), .D(n1754), 
        .Q(readOutBus[583]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_104_ ( .G(n2006), .D(n1756), 
        .Q(readOutBus[584]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_105_ ( .G(n2006), .D(n1758), 
        .Q(readOutBus[585]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_106_ ( .G(n2006), .D(n1760), 
        .Q(readOutBus[586]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_107_ ( .G(n2006), .D(n1762), 
        .Q(readOutBus[587]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_112_ ( .G(n2004), .D(n1772), 
        .Q(readOutBus[592]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_113_ ( .G(n2004), .D(n1774), 
        .Q(readOutBus[593]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_114_ ( .G(n2004), .D(n1776), 
        .Q(readOutBus[594]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_115_ ( .G(n2004), .D(n1778), 
        .Q(readOutBus[595]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_156_ ( .G(n1994), .D(n1860), 
        .Q(readOutBus[636]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_157_ ( .G(n1994), .D(n1862), 
        .Q(readOutBus[637]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_158_ ( .G(n1994), .D(n1864), 
        .Q(readOutBus[638]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_159_ ( .G(n1994), .D(n1866), 
        .Q(readOutBus[639]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_24_ ( .G(n2102), .D(n1596), 
        .Q(readOutBus[824]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_25_ ( .G(n2102), .D(n1598), 
        .Q(readOutBus[825]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_26_ ( .G(n2102), .D(n1600), 
        .Q(readOutBus[826]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_27_ ( .G(n2102), .D(n1602), 
        .Q(readOutBus[827]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_28_ ( .G(n2101), .D(n1604), 
        .Q(readOutBus[828]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_29_ ( .G(n2101), .D(n1606), 
        .Q(readOutBus[829]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_30_ ( .G(n2101), .D(n1608), 
        .Q(readOutBus[830]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_31_ ( .G(n2101), .D(n1610), 
        .Q(readOutBus[831]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_32_ ( .G(n2100), .D(n1612), 
        .Q(readOutBus[832]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_33_ ( .G(n2100), .D(n1614), 
        .Q(readOutBus[833]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_34_ ( .G(n2100), .D(n1616), 
        .Q(readOutBus[834]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_35_ ( .G(n2100), .D(n1618), 
        .Q(readOutBus[835]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_40_ ( .G(n2098), .D(n1628), 
        .Q(readOutBus[840]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_41_ ( .G(n2098), .D(n1630), 
        .Q(readOutBus[841]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_42_ ( .G(n2098), .D(n1632), 
        .Q(readOutBus[842]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_43_ ( .G(n2098), .D(n1634), 
        .Q(readOutBus[843]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_48_ ( .G(n2096), .D(n1644), 
        .Q(readOutBus[848]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_49_ ( .G(n2096), .D(n1646), 
        .Q(readOutBus[849]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_50_ ( .G(n2096), .D(n1648), 
        .Q(readOutBus[850]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_51_ ( .G(n2096), .D(n1650), 
        .Q(readOutBus[851]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_52_ ( .G(n2095), .D(n1652), 
        .Q(readOutBus[852]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_53_ ( .G(n2095), .D(n1654), 
        .Q(readOutBus[853]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_54_ ( .G(n2095), .D(n1656), 
        .Q(readOutBus[854]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_55_ ( .G(n2095), .D(n1658), 
        .Q(readOutBus[855]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_56_ ( .G(n2094), .D(n1660), 
        .Q(readOutBus[856]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_57_ ( .G(n2094), .D(n1662), 
        .Q(readOutBus[857]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_58_ ( .G(n2094), .D(n1664), 
        .Q(readOutBus[858]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_59_ ( .G(n2094), .D(n1666), 
        .Q(readOutBus[859]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_60_ ( .G(n2093), .D(n1668), 
        .Q(readOutBus[860]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_61_ ( .G(n2093), .D(n1670), 
        .Q(readOutBus[861]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_62_ ( .G(n2093), .D(n1672), 
        .Q(readOutBus[862]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_63_ ( .G(n2093), .D(n1674), 
        .Q(readOutBus[863]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_64_ ( .G(n2092), .D(n1676), 
        .Q(readOutBus[864]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_65_ ( .G(n2092), .D(n1678), 
        .Q(readOutBus[865]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_66_ ( .G(n2092), .D(n1680), 
        .Q(readOutBus[866]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_67_ ( .G(n2092), .D(n1682), 
        .Q(readOutBus[867]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_68_ ( .G(n2091), .D(n1684), 
        .Q(readOutBus[868]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_69_ ( .G(n2091), .D(n1686), 
        .Q(readOutBus[869]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_70_ ( .G(n2091), .D(n1688), 
        .Q(readOutBus[870]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_71_ ( .G(n2091), .D(n1690), 
        .Q(readOutBus[871]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_72_ ( .G(n2090), .D(n1692), 
        .Q(readOutBus[872]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_73_ ( .G(n2090), .D(n1694), 
        .Q(readOutBus[873]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_74_ ( .G(n2090), .D(n1696), 
        .Q(readOutBus[874]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_75_ ( .G(n2090), .D(n1698), 
        .Q(readOutBus[875]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_96_ ( .G(n2084), .D(n1740), 
        .Q(readOutBus[896]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_97_ ( .G(n2084), .D(n1742), 
        .Q(readOutBus[897]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_98_ ( .G(n2084), .D(n1744), 
        .Q(readOutBus[898]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_99_ ( .G(n2084), .D(n1746), 
        .Q(readOutBus[899]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_100_ ( .G(n2083), .D(n1748), 
        .Q(readOutBus[900]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_101_ ( .G(n2083), .D(n1750), 
        .Q(readOutBus[901]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_102_ ( .G(n2083), .D(n1752), 
        .Q(readOutBus[902]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_103_ ( .G(n2083), .D(n1754), 
        .Q(readOutBus[903]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_104_ ( .G(n2082), .D(n1756), 
        .Q(readOutBus[904]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_105_ ( .G(n2082), .D(n1758), 
        .Q(readOutBus[905]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_106_ ( .G(n2082), .D(n1760), 
        .Q(readOutBus[906]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_107_ ( .G(n2082), .D(n1762), 
        .Q(readOutBus[907]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_112_ ( .G(n2080), .D(n1772), 
        .Q(readOutBus[912]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_113_ ( .G(n2080), .D(n1774), 
        .Q(readOutBus[913]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_114_ ( .G(n2080), .D(n1776), 
        .Q(readOutBus[914]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_115_ ( .G(n2080), .D(n1778), 
        .Q(readOutBus[915]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_136_ ( .G(n2075), .D(n1820), 
        .Q(readOutBus[936]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_137_ ( .G(n2075), .D(n1822), 
        .Q(readOutBus[937]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_138_ ( .G(n2075), .D(n1824), 
        .Q(readOutBus[938]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_139_ ( .G(n2075), .D(n1826), 
        .Q(readOutBus[939]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_140_ ( .G(n2074), .D(n1828), 
        .Q(readOutBus[940]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_141_ ( .G(n2074), .D(n1830), 
        .Q(readOutBus[941]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_142_ ( .G(n2074), .D(n1832), 
        .Q(readOutBus[942]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_143_ ( .G(n2074), .D(n1834), 
        .Q(readOutBus[943]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_144_ ( .G(n2073), .D(n1836), 
        .Q(readOutBus[944]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_145_ ( .G(n2073), .D(n1838), 
        .Q(readOutBus[945]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_146_ ( .G(n2073), .D(n1840), 
        .Q(readOutBus[946]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_147_ ( .G(n2073), .D(n1842), 
        .Q(readOutBus[947]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_156_ ( .G(n2070), .D(n1860), 
        .Q(readOutBus[956]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_157_ ( .G(n2070), .D(n1862), 
        .Q(readOutBus[957]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_158_ ( .G(n2070), .D(n1864), 
        .Q(readOutBus[958]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_159_ ( .G(n2070), .D(n1866), 
        .Q(readOutBus[959]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_0_ ( .G(n1955), .D(n1548), 
        .Q(readOutBus[160]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_1_ ( .G(n1955), .D(n1550), 
        .Q(readOutBus[161]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_2_ ( .G(n1955), .D(n1552), 
        .Q(readOutBus[162]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_3_ ( .G(n1955), .D(n1554), 
        .Q(readOutBus[163]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_8_ ( .G(n1954), .D(n1564), 
        .Q(readOutBus[168]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_9_ ( .G(n1954), .D(n1566), 
        .Q(readOutBus[169]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_10_ ( .G(n1954), .D(n1568), 
        .Q(readOutBus[170]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_11_ ( .G(n1954), .D(n1570), 
        .Q(readOutBus[171]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_36_ ( .G(n1947), .D(n1620), 
        .Q(readOutBus[196]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_37_ ( .G(n1947), .D(n1622), 
        .Q(readOutBus[197]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_38_ ( .G(n1947), .D(n1624), 
        .Q(readOutBus[198]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_39_ ( .G(n1947), .D(n1626), 
        .Q(readOutBus[199]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_80_ ( .G(n1936), .D(n1708), 
        .Q(readOutBus[240]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_81_ ( .G(n1936), .D(n1710), 
        .Q(readOutBus[241]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_82_ ( .G(n1936), .D(n1712), 
        .Q(readOutBus[242]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_83_ ( .G(n1936), .D(n1714), 
        .Q(readOutBus[243]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_108_ ( .G(n1929), .D(n1764), 
        .Q(readOutBus[268]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_109_ ( .G(n1929), .D(n1766), 
        .Q(readOutBus[269]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_110_ ( .G(n1929), .D(n1768), 
        .Q(readOutBus[270]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_111_ ( .G(n1929), .D(n1770), 
        .Q(readOutBus[271]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_116_ ( .G(n1927), .D(n1780), 
        .Q(readOutBus[276]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_117_ ( .G(n1927), .D(n1782), 
        .Q(readOutBus[277]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_118_ ( .G(n1927), .D(n1784), 
        .Q(readOutBus[278]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_119_ ( .G(n1927), .D(n1786), 
        .Q(readOutBus[279]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_148_ ( .G(n1920), .D(n1844), 
        .Q(readOutBus[308]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_149_ ( .G(n1920), .D(n1846), 
        .Q(readOutBus[309]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_150_ ( .G(n1920), .D(n1848), 
        .Q(readOutBus[310]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_151_ ( .G(n1920), .D(n1850), 
        .Q(readOutBus[311]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_0_ ( .G(n2031), .D(n1548), 
        .Q(readOutBus[480]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_1_ ( .G(n2031), .D(n1550), 
        .Q(readOutBus[481]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_2_ ( .G(n2031), .D(n1552), 
        .Q(readOutBus[482]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_3_ ( .G(n2031), .D(n1554), 
        .Q(readOutBus[483]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_8_ ( .G(n2030), .D(n1564), 
        .Q(readOutBus[488]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_9_ ( .G(n2030), .D(n1566), 
        .Q(readOutBus[489]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_10_ ( .G(n2030), .D(n1568), 
        .Q(readOutBus[490]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_11_ ( .G(n2030), .D(n1570), 
        .Q(readOutBus[491]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_36_ ( .G(n2023), .D(n1620), 
        .Q(readOutBus[516]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_37_ ( .G(n2023), .D(n1622), 
        .Q(readOutBus[517]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_38_ ( .G(n2023), .D(n1624), 
        .Q(readOutBus[518]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_39_ ( .G(n2023), .D(n1626), 
        .Q(readOutBus[519]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_80_ ( .G(n2012), .D(n1708), 
        .Q(readOutBus[560]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_81_ ( .G(n2012), .D(n1710), 
        .Q(readOutBus[561]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_82_ ( .G(n2012), .D(n1712), 
        .Q(readOutBus[562]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_83_ ( .G(n2012), .D(n1714), 
        .Q(readOutBus[563]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_108_ ( .G(n2005), .D(n1764), 
        .Q(readOutBus[588]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_109_ ( .G(n2005), .D(n1766), 
        .Q(readOutBus[589]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_110_ ( .G(n2005), .D(n1768), 
        .Q(readOutBus[590]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_111_ ( .G(n2005), .D(n1770), 
        .Q(readOutBus[591]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_116_ ( .G(n2003), .D(n1780), 
        .Q(readOutBus[596]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_117_ ( .G(n2003), .D(n1782), 
        .Q(readOutBus[597]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_118_ ( .G(n2003), .D(n1784), 
        .Q(readOutBus[598]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_119_ ( .G(n2003), .D(n1786), 
        .Q(readOutBus[599]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_148_ ( .G(n1996), .D(n1844), 
        .Q(readOutBus[628]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_149_ ( .G(n1996), .D(n1846), 
        .Q(readOutBus[629]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_150_ ( .G(n1996), .D(n1848), 
        .Q(readOutBus[630]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_151_ ( .G(n1996), .D(n1850), 
        .Q(readOutBus[631]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_0_ ( .G(n2107), .D(n1548), 
        .Q(readOutBus[800]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_1_ ( .G(n2107), .D(n1550), 
        .Q(readOutBus[801]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_2_ ( .G(n2107), .D(n1552), 
        .Q(readOutBus[802]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_3_ ( .G(n2107), .D(n1554), 
        .Q(readOutBus[803]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_8_ ( .G(n2106), .D(n1564), 
        .Q(readOutBus[808]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_9_ ( .G(n2106), .D(n1566), 
        .Q(readOutBus[809]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_10_ ( .G(n2106), .D(n1568), 
        .Q(readOutBus[810]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_11_ ( .G(n2106), .D(n1570), 
        .Q(readOutBus[811]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_132_ ( .G(n2076), .D(n1812), 
        .Q(readOutBus[932]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_133_ ( .G(n2076), .D(n1814), 
        .Q(readOutBus[933]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_134_ ( .G(n2076), .D(n1816), 
        .Q(readOutBus[934]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_135_ ( .G(n2076), .D(n1818), 
        .Q(readOutBus[935]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_5_ ( .G(n1870), .D(n1558), 
        .Q(readOutBus[165]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_7_ ( .G(n1870), .D(n1562), 
        .Q(readOutBus[167]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_5_ ( .G(n1874), .D(n1558), 
        .Q(readOutBus[485]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_7_ ( .G(n1874), .D(n1562), 
        .Q(readOutBus[487]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_5_ ( .G(n1878), .D(n1558), 
        .Q(readOutBus[805]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_7_ ( .G(n1878), .D(n1562), 
        .Q(readOutBus[807]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_36_ ( .G(n2099), .D(n1620), 
        .Q(readOutBus[836]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_37_ ( .G(n2099), .D(n1622), 
        .Q(readOutBus[837]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_38_ ( .G(n2099), .D(n1624), 
        .Q(readOutBus[838]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_39_ ( .G(n2099), .D(n1626), 
        .Q(readOutBus[839]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_80_ ( .G(n2088), .D(n1708), 
        .Q(readOutBus[880]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_81_ ( .G(n2088), .D(n1710), 
        .Q(readOutBus[881]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_82_ ( .G(n2088), .D(n1712), 
        .Q(readOutBus[882]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_83_ ( .G(n2088), .D(n1714), 
        .Q(readOutBus[883]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_108_ ( .G(n2081), .D(n1764), 
        .Q(readOutBus[908]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_109_ ( .G(n2081), .D(n1766), 
        .Q(readOutBus[909]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_110_ ( .G(n2081), .D(n1768), 
        .Q(readOutBus[910]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_111_ ( .G(n2081), .D(n1770), 
        .Q(readOutBus[911]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_116_ ( .G(n2079), .D(n1780), 
        .Q(readOutBus[916]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_117_ ( .G(n2079), .D(n1782), 
        .Q(readOutBus[917]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_118_ ( .G(n2079), .D(n1784), 
        .Q(readOutBus[918]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_119_ ( .G(n2079), .D(n1786), 
        .Q(readOutBus[919]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_148_ ( .G(n2072), .D(n1844), 
        .Q(readOutBus[948]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_149_ ( .G(n2072), .D(n1846), 
        .Q(readOutBus[949]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_150_ ( .G(n2072), .D(n1848), 
        .Q(readOutBus[950]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_151_ ( .G(n2072), .D(n1850), 
        .Q(readOutBus[951]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_152_ ( .G(n2071), .D(n1852), 
        .Q(readOutBus[952]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_153_ ( .G(n2071), .D(n1854), 
        .Q(readOutBus[953]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_154_ ( .G(n2071), .D(n1856), 
        .Q(readOutBus[954]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_155_ ( .G(n2071), .D(n1858), 
        .Q(readOutBus[955]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_12_ ( .G(n1953), .D(n1572), 
        .Q(readOutBus[172]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_13_ ( .G(n1953), .D(n1574), 
        .Q(readOutBus[173]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_14_ ( .G(n1953), .D(n1576), 
        .Q(readOutBus[174]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_15_ ( .G(n1953), .D(n1578), 
        .Q(readOutBus[175]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_16_ ( .G(n1952), .D(n1580), 
        .Q(readOutBus[176]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_17_ ( .G(n1952), .D(n1582), 
        .Q(readOutBus[177]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_18_ ( .G(n1952), .D(n1584), 
        .Q(readOutBus[178]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_19_ ( .G(n1952), .D(n1586), 
        .Q(readOutBus[179]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_20_ ( .G(n1951), .D(n1588), 
        .Q(readOutBus[180]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_21_ ( .G(n1951), .D(n1590), 
        .Q(readOutBus[181]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_22_ ( .G(n1951), .D(n1592), 
        .Q(readOutBus[182]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_23_ ( .G(n1951), .D(n1594), 
        .Q(readOutBus[183]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_48_ ( .G(n1944), .D(n1644), 
        .Q(readOutBus[208]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_49_ ( .G(n1944), .D(n1646), 
        .Q(readOutBus[209]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_50_ ( .G(n1944), .D(n1648), 
        .Q(readOutBus[210]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_51_ ( .G(n1944), .D(n1650), 
        .Q(readOutBus[211]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_52_ ( .G(n1943), .D(n1652), 
        .Q(readOutBus[212]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_53_ ( .G(n1943), .D(n1654), 
        .Q(readOutBus[213]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_54_ ( .G(n1943), .D(n1656), 
        .Q(readOutBus[214]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_55_ ( .G(n1943), .D(n1658), 
        .Q(readOutBus[215]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_56_ ( .G(n1942), .D(n1660), 
        .Q(readOutBus[216]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_57_ ( .G(n1942), .D(n1662), 
        .Q(readOutBus[217]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_58_ ( .G(n1942), .D(n1664), 
        .Q(readOutBus[218]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_59_ ( .G(n1942), .D(n1666), 
        .Q(readOutBus[219]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_12_ ( .G(n2029), .D(n1572), 
        .Q(readOutBus[492]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_13_ ( .G(n2029), .D(n1574), 
        .Q(readOutBus[493]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_14_ ( .G(n2029), .D(n1576), 
        .Q(readOutBus[494]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_15_ ( .G(n2029), .D(n1578), 
        .Q(readOutBus[495]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_16_ ( .G(n2028), .D(n1580), 
        .Q(readOutBus[496]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_17_ ( .G(n2028), .D(n1582), 
        .Q(readOutBus[497]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_18_ ( .G(n2028), .D(n1584), 
        .Q(readOutBus[498]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_19_ ( .G(n2028), .D(n1586), 
        .Q(readOutBus[499]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_20_ ( .G(n2027), .D(n1588), 
        .Q(readOutBus[500]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_21_ ( .G(n2027), .D(n1590), 
        .Q(readOutBus[501]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_22_ ( .G(n2027), .D(n1592), 
        .Q(readOutBus[502]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_23_ ( .G(n2027), .D(n1594), 
        .Q(readOutBus[503]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_48_ ( .G(n2020), .D(n1644), 
        .Q(readOutBus[528]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_49_ ( .G(n2020), .D(n1646), 
        .Q(readOutBus[529]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_50_ ( .G(n2020), .D(n1648), 
        .Q(readOutBus[530]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_51_ ( .G(n2020), .D(n1650), 
        .Q(readOutBus[531]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_52_ ( .G(n2019), .D(n1652), 
        .Q(readOutBus[532]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_53_ ( .G(n2019), .D(n1654), 
        .Q(readOutBus[533]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_54_ ( .G(n2019), .D(n1656), 
        .Q(readOutBus[534]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_55_ ( .G(n2019), .D(n1658), 
        .Q(readOutBus[535]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_56_ ( .G(n2018), .D(n1660), 
        .Q(readOutBus[536]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_57_ ( .G(n2018), .D(n1662), 
        .Q(readOutBus[537]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_58_ ( .G(n2018), .D(n1664), 
        .Q(readOutBus[538]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_59_ ( .G(n2018), .D(n1666), 
        .Q(readOutBus[539]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_12_ ( .G(n2105), .D(n1572), 
        .Q(readOutBus[812]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_13_ ( .G(n2105), .D(n1574), 
        .Q(readOutBus[813]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_14_ ( .G(n2105), .D(n1576), 
        .Q(readOutBus[814]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_15_ ( .G(n2105), .D(n1578), 
        .Q(readOutBus[815]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_16_ ( .G(n2104), .D(n1580), 
        .Q(readOutBus[816]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_17_ ( .G(n2104), .D(n1582), 
        .Q(readOutBus[817]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_18_ ( .G(n2104), .D(n1584), 
        .Q(readOutBus[818]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_19_ ( .G(n2104), .D(n1586), 
        .Q(readOutBus[819]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_20_ ( .G(n2103), .D(n1588), 
        .Q(readOutBus[820]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_21_ ( .G(n2103), .D(n1590), 
        .Q(readOutBus[821]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_22_ ( .G(n2103), .D(n1592), 
        .Q(readOutBus[822]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_23_ ( .G(n2103), .D(n1594), 
        .Q(readOutBus[823]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_4_ ( .G(n1871), .D(n1556), 
        .Q(readOutBus[164]) );
  TLATXLTS Generate_Node_Banks_1__NB_readOut_reg_6_ ( .G(n1871), .D(n1560), 
        .Q(readOutBus[166]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_4_ ( .G(n1875), .D(n1556), 
        .Q(readOutBus[484]) );
  TLATXLTS Generate_Node_Banks_3__NB_readOut_reg_6_ ( .G(n1875), .D(n1560), 
        .Q(readOutBus[486]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_4_ ( .G(n1879), .D(n1556), 
        .Q(readOutBus[804]) );
  TLATXLTS Generate_Node_Banks_5__NB_readOut_reg_6_ ( .G(n1879), .D(n1560), 
        .Q(readOutBus[806]) );
  INVX2TS U664 ( .A(writeIn[0]), .Y(n496) );
  INVX2TS U665 ( .A(n496), .Y(n1548) );
  INVX2TS U666 ( .A(n496), .Y(n1549) );
  INVX2TS U667 ( .A(writeIn[1]), .Y(n497) );
  INVX2TS U668 ( .A(n497), .Y(n1550) );
  INVX2TS U669 ( .A(n497), .Y(n1551) );
  INVX2TS U670 ( .A(writeIn[2]), .Y(n498) );
  INVX2TS U671 ( .A(n498), .Y(n1552) );
  INVX2TS U672 ( .A(n498), .Y(n1553) );
  INVX2TS U673 ( .A(writeIn[3]), .Y(n499) );
  INVX2TS U674 ( .A(n499), .Y(n1554) );
  INVX2TS U675 ( .A(n499), .Y(n1555) );
  INVX2TS U676 ( .A(writeIn[4]), .Y(n500) );
  INVX2TS U677 ( .A(n500), .Y(n1556) );
  INVX2TS U678 ( .A(n500), .Y(n1557) );
  INVX2TS U679 ( .A(writeIn[5]), .Y(n501) );
  INVX2TS U680 ( .A(n501), .Y(n1558) );
  INVX2TS U681 ( .A(n501), .Y(n1559) );
  INVX2TS U682 ( .A(writeIn[6]), .Y(n502) );
  INVX2TS U683 ( .A(n502), .Y(n1560) );
  INVX2TS U684 ( .A(n502), .Y(n1561) );
  INVX2TS U685 ( .A(writeIn[7]), .Y(n503) );
  INVX2TS U686 ( .A(n503), .Y(n1562) );
  INVX2TS U687 ( .A(n503), .Y(n1563) );
  INVX2TS U688 ( .A(writeIn[8]), .Y(n504) );
  INVX2TS U689 ( .A(n504), .Y(n1564) );
  INVX2TS U690 ( .A(n504), .Y(n1565) );
  INVX2TS U691 ( .A(writeIn[9]), .Y(n505) );
  INVX2TS U692 ( .A(n505), .Y(n1566) );
  INVX2TS U693 ( .A(n505), .Y(n1567) );
  INVX2TS U694 ( .A(writeIn[10]), .Y(n506) );
  INVX2TS U695 ( .A(n506), .Y(n1568) );
  INVX2TS U696 ( .A(n506), .Y(n1569) );
  INVX2TS U697 ( .A(writeIn[11]), .Y(n507) );
  INVX2TS U698 ( .A(n507), .Y(n1570) );
  INVX2TS U699 ( .A(n507), .Y(n1571) );
  INVX2TS U700 ( .A(writeIn[12]), .Y(n508) );
  INVX2TS U701 ( .A(n508), .Y(n1572) );
  INVX2TS U702 ( .A(n508), .Y(n1573) );
  INVX2TS U703 ( .A(writeIn[13]), .Y(n509) );
  INVX2TS U704 ( .A(n509), .Y(n1574) );
  INVX2TS U705 ( .A(n509), .Y(n1575) );
  INVX2TS U706 ( .A(writeIn[14]), .Y(n510) );
  INVX2TS U707 ( .A(n510), .Y(n1576) );
  INVX2TS U708 ( .A(n510), .Y(n1577) );
  INVX2TS U709 ( .A(writeIn[15]), .Y(n511) );
  INVX2TS U710 ( .A(n511), .Y(n1578) );
  INVX2TS U711 ( .A(n511), .Y(n1579) );
  INVX2TS U712 ( .A(writeIn[16]), .Y(n512) );
  INVX2TS U713 ( .A(n512), .Y(n1580) );
  INVX2TS U714 ( .A(n512), .Y(n1581) );
  INVX2TS U715 ( .A(writeIn[17]), .Y(n513) );
  INVX2TS U716 ( .A(n513), .Y(n1582) );
  INVX2TS U717 ( .A(n513), .Y(n1583) );
  INVX2TS U718 ( .A(writeIn[18]), .Y(n514) );
  INVX2TS U719 ( .A(n514), .Y(n1584) );
  INVX2TS U720 ( .A(n514), .Y(n1585) );
  INVX2TS U721 ( .A(writeIn[19]), .Y(n515) );
  INVX2TS U722 ( .A(n515), .Y(n1586) );
  INVX2TS U723 ( .A(n515), .Y(n1587) );
  INVX2TS U724 ( .A(writeIn[20]), .Y(n516) );
  INVX2TS U725 ( .A(n516), .Y(n1588) );
  INVX2TS U726 ( .A(n516), .Y(n1589) );
  INVX2TS U727 ( .A(writeIn[21]), .Y(n517) );
  INVX2TS U728 ( .A(n517), .Y(n1590) );
  INVX2TS U729 ( .A(n517), .Y(n1591) );
  INVX2TS U730 ( .A(writeIn[22]), .Y(n518) );
  INVX2TS U731 ( .A(n518), .Y(n1592) );
  INVX2TS U732 ( .A(n518), .Y(n1593) );
  INVX2TS U733 ( .A(writeIn[23]), .Y(n519) );
  INVX2TS U734 ( .A(n519), .Y(n1594) );
  INVX2TS U735 ( .A(n519), .Y(n1595) );
  INVX2TS U736 ( .A(writeIn[24]), .Y(n520) );
  INVX2TS U737 ( .A(n520), .Y(n1596) );
  INVX2TS U738 ( .A(n520), .Y(n1597) );
  INVX2TS U739 ( .A(writeIn[25]), .Y(n521) );
  INVX2TS U740 ( .A(n521), .Y(n1598) );
  INVX2TS U741 ( .A(n521), .Y(n1599) );
  INVX2TS U742 ( .A(writeIn[26]), .Y(n522) );
  INVX2TS U743 ( .A(n522), .Y(n1600) );
  INVX2TS U744 ( .A(n522), .Y(n1601) );
  INVX2TS U745 ( .A(writeIn[27]), .Y(n523) );
  INVX2TS U746 ( .A(n523), .Y(n1602) );
  INVX2TS U747 ( .A(n523), .Y(n1603) );
  INVX2TS U748 ( .A(writeIn[28]), .Y(n524) );
  INVX2TS U749 ( .A(n524), .Y(n1604) );
  INVX2TS U750 ( .A(n524), .Y(n1605) );
  INVX2TS U751 ( .A(writeIn[29]), .Y(n525) );
  INVX2TS U752 ( .A(n525), .Y(n1606) );
  INVX2TS U753 ( .A(n525), .Y(n1607) );
  INVX2TS U754 ( .A(writeIn[30]), .Y(n526) );
  INVX2TS U755 ( .A(n526), .Y(n1608) );
  INVX2TS U756 ( .A(n526), .Y(n1609) );
  INVX2TS U757 ( .A(writeIn[31]), .Y(n527) );
  INVX2TS U758 ( .A(n527), .Y(n1610) );
  INVX2TS U759 ( .A(n527), .Y(n1611) );
  INVX2TS U760 ( .A(writeIn[32]), .Y(n528) );
  INVX2TS U761 ( .A(n528), .Y(n1612) );
  INVX2TS U762 ( .A(n528), .Y(n1613) );
  INVX2TS U763 ( .A(writeIn[33]), .Y(n529) );
  INVX2TS U764 ( .A(n529), .Y(n1614) );
  INVX2TS U765 ( .A(n529), .Y(n1615) );
  INVX2TS U766 ( .A(writeIn[34]), .Y(n530) );
  INVX2TS U767 ( .A(n530), .Y(n1616) );
  INVX2TS U768 ( .A(n530), .Y(n1617) );
  INVX2TS U769 ( .A(writeIn[35]), .Y(n531) );
  INVX2TS U770 ( .A(n531), .Y(n1618) );
  INVX2TS U771 ( .A(n531), .Y(n1619) );
  INVX2TS U772 ( .A(writeIn[36]), .Y(n532) );
  INVX2TS U773 ( .A(n532), .Y(n1620) );
  INVX2TS U774 ( .A(n532), .Y(n1621) );
  INVX2TS U775 ( .A(writeIn[37]), .Y(n533) );
  INVX2TS U776 ( .A(n533), .Y(n1622) );
  INVX2TS U777 ( .A(n533), .Y(n1623) );
  INVX2TS U778 ( .A(writeIn[38]), .Y(n534) );
  INVX2TS U779 ( .A(n534), .Y(n1624) );
  INVX2TS U780 ( .A(n534), .Y(n1625) );
  INVX2TS U781 ( .A(writeIn[39]), .Y(n535) );
  INVX2TS U782 ( .A(n535), .Y(n1626) );
  INVX2TS U783 ( .A(n535), .Y(n1627) );
  INVX2TS U784 ( .A(writeIn[40]), .Y(n536) );
  INVX2TS U785 ( .A(n536), .Y(n1628) );
  INVX2TS U786 ( .A(n536), .Y(n1629) );
  INVX2TS U787 ( .A(writeIn[41]), .Y(n537) );
  INVX2TS U788 ( .A(n537), .Y(n1630) );
  INVX2TS U789 ( .A(n537), .Y(n1631) );
  INVX2TS U790 ( .A(writeIn[42]), .Y(n538) );
  INVX2TS U791 ( .A(n538), .Y(n1632) );
  INVX2TS U792 ( .A(n538), .Y(n1633) );
  INVX2TS U793 ( .A(writeIn[43]), .Y(n539) );
  INVX2TS U794 ( .A(n539), .Y(n1634) );
  INVX2TS U795 ( .A(n539), .Y(n1635) );
  INVX2TS U796 ( .A(writeIn[44]), .Y(n540) );
  INVX2TS U797 ( .A(n540), .Y(n1636) );
  INVX2TS U798 ( .A(n540), .Y(n1637) );
  INVX2TS U799 ( .A(writeIn[45]), .Y(n541) );
  INVX2TS U800 ( .A(n541), .Y(n1638) );
  INVX2TS U801 ( .A(n541), .Y(n1639) );
  INVX2TS U802 ( .A(writeIn[46]), .Y(n542) );
  INVX2TS U803 ( .A(n542), .Y(n1640) );
  INVX2TS U804 ( .A(n542), .Y(n1641) );
  INVX2TS U805 ( .A(writeIn[47]), .Y(n543) );
  INVX2TS U806 ( .A(n543), .Y(n1642) );
  INVX2TS U807 ( .A(n543), .Y(n1643) );
  INVX2TS U808 ( .A(writeIn[48]), .Y(n544) );
  INVX2TS U809 ( .A(n544), .Y(n1644) );
  INVX2TS U810 ( .A(n544), .Y(n1645) );
  INVX2TS U811 ( .A(writeIn[49]), .Y(n545) );
  INVX2TS U812 ( .A(n545), .Y(n1646) );
  INVX2TS U813 ( .A(n545), .Y(n1647) );
  INVX2TS U814 ( .A(writeIn[50]), .Y(n546) );
  INVX2TS U815 ( .A(n546), .Y(n1648) );
  INVX2TS U816 ( .A(n546), .Y(n1649) );
  INVX2TS U817 ( .A(writeIn[51]), .Y(n547) );
  INVX2TS U818 ( .A(n547), .Y(n1650) );
  INVX2TS U819 ( .A(n547), .Y(n1651) );
  INVX2TS U820 ( .A(writeIn[52]), .Y(n548) );
  INVX2TS U821 ( .A(n548), .Y(n1652) );
  INVX2TS U822 ( .A(n548), .Y(n1653) );
  INVX2TS U823 ( .A(writeIn[53]), .Y(n549) );
  INVX2TS U824 ( .A(n549), .Y(n1654) );
  INVX2TS U825 ( .A(n549), .Y(n1655) );
  INVX2TS U826 ( .A(writeIn[54]), .Y(n550) );
  INVX2TS U827 ( .A(n550), .Y(n1656) );
  INVX2TS U828 ( .A(n550), .Y(n1657) );
  INVX2TS U829 ( .A(writeIn[55]), .Y(n551) );
  INVX2TS U830 ( .A(n551), .Y(n1658) );
  INVX2TS U831 ( .A(n551), .Y(n1659) );
  INVX2TS U832 ( .A(writeIn[56]), .Y(n552) );
  INVX2TS U833 ( .A(n552), .Y(n1660) );
  INVX2TS U834 ( .A(n552), .Y(n1661) );
  INVX2TS U835 ( .A(writeIn[57]), .Y(n553) );
  INVX2TS U836 ( .A(n553), .Y(n1662) );
  INVX2TS U837 ( .A(n553), .Y(n1663) );
  INVX2TS U838 ( .A(writeIn[58]), .Y(n554) );
  INVX2TS U839 ( .A(n554), .Y(n1664) );
  INVX2TS U840 ( .A(n554), .Y(n1665) );
  INVX2TS U841 ( .A(writeIn[59]), .Y(n555) );
  INVX2TS U842 ( .A(n555), .Y(n1666) );
  INVX2TS U843 ( .A(n555), .Y(n1667) );
  INVX2TS U844 ( .A(writeIn[60]), .Y(n556) );
  INVX2TS U845 ( .A(n556), .Y(n1668) );
  INVX2TS U846 ( .A(n556), .Y(n1669) );
  INVX2TS U847 ( .A(writeIn[61]), .Y(n557) );
  INVX2TS U848 ( .A(n557), .Y(n1670) );
  INVX2TS U849 ( .A(n557), .Y(n1671) );
  INVX2TS U850 ( .A(writeIn[62]), .Y(n558) );
  INVX2TS U851 ( .A(n558), .Y(n1672) );
  INVX2TS U852 ( .A(n558), .Y(n1673) );
  INVX2TS U853 ( .A(writeIn[63]), .Y(n559) );
  INVX2TS U854 ( .A(n559), .Y(n1674) );
  INVX2TS U855 ( .A(n559), .Y(n1675) );
  INVX2TS U856 ( .A(writeIn[64]), .Y(n560) );
  INVX2TS U857 ( .A(n560), .Y(n1676) );
  INVX2TS U858 ( .A(n560), .Y(n1677) );
  INVX2TS U859 ( .A(writeIn[65]), .Y(n561) );
  INVX2TS U860 ( .A(n561), .Y(n1678) );
  INVX2TS U861 ( .A(n561), .Y(n1679) );
  INVX2TS U862 ( .A(writeIn[66]), .Y(n562) );
  INVX2TS U863 ( .A(n562), .Y(n1680) );
  INVX2TS U864 ( .A(n562), .Y(n1681) );
  INVX2TS U865 ( .A(writeIn[67]), .Y(n563) );
  INVX2TS U866 ( .A(n563), .Y(n1682) );
  INVX2TS U867 ( .A(n563), .Y(n1683) );
  INVX2TS U868 ( .A(writeIn[68]), .Y(n564) );
  INVX2TS U869 ( .A(n564), .Y(n1684) );
  INVX2TS U870 ( .A(n564), .Y(n1685) );
  INVX2TS U871 ( .A(writeIn[69]), .Y(n565) );
  INVX2TS U872 ( .A(n565), .Y(n1686) );
  INVX2TS U873 ( .A(n565), .Y(n1687) );
  INVX2TS U874 ( .A(writeIn[70]), .Y(n566) );
  INVX2TS U875 ( .A(n566), .Y(n1688) );
  INVX2TS U876 ( .A(n566), .Y(n1689) );
  INVX2TS U877 ( .A(writeIn[71]), .Y(n567) );
  INVX2TS U878 ( .A(n567), .Y(n1690) );
  INVX2TS U879 ( .A(n567), .Y(n1691) );
  INVX2TS U880 ( .A(writeIn[72]), .Y(n568) );
  INVX2TS U881 ( .A(n568), .Y(n1692) );
  INVX2TS U882 ( .A(n568), .Y(n1693) );
  INVX2TS U883 ( .A(writeIn[73]), .Y(n569) );
  INVX2TS U884 ( .A(n569), .Y(n1694) );
  INVX2TS U885 ( .A(n569), .Y(n1695) );
  INVX2TS U886 ( .A(writeIn[74]), .Y(n570) );
  INVX2TS U887 ( .A(n570), .Y(n1696) );
  INVX2TS U888 ( .A(n570), .Y(n1697) );
  INVX2TS U889 ( .A(writeIn[75]), .Y(n571) );
  INVX2TS U890 ( .A(n571), .Y(n1698) );
  INVX2TS U891 ( .A(n571), .Y(n1699) );
  INVX2TS U892 ( .A(writeIn[76]), .Y(n572) );
  INVX2TS U893 ( .A(n572), .Y(n1700) );
  INVX2TS U894 ( .A(n572), .Y(n1701) );
  INVX2TS U895 ( .A(writeIn[77]), .Y(n573) );
  INVX2TS U896 ( .A(n573), .Y(n1702) );
  INVX2TS U897 ( .A(n573), .Y(n1703) );
  INVX2TS U898 ( .A(writeIn[78]), .Y(n574) );
  INVX2TS U899 ( .A(n574), .Y(n1704) );
  INVX2TS U900 ( .A(n574), .Y(n1705) );
  INVX2TS U901 ( .A(writeIn[79]), .Y(n575) );
  INVX2TS U902 ( .A(n575), .Y(n1706) );
  INVX2TS U903 ( .A(n575), .Y(n1707) );
  INVX2TS U904 ( .A(writeIn[80]), .Y(n576) );
  INVX2TS U905 ( .A(n576), .Y(n1708) );
  INVX2TS U906 ( .A(n576), .Y(n1709) );
  INVX2TS U907 ( .A(writeIn[81]), .Y(n577) );
  INVX2TS U908 ( .A(n577), .Y(n1710) );
  INVX2TS U909 ( .A(n577), .Y(n1711) );
  INVX2TS U910 ( .A(writeIn[82]), .Y(n578) );
  INVX2TS U911 ( .A(n578), .Y(n1712) );
  INVX2TS U912 ( .A(n578), .Y(n1713) );
  INVX2TS U913 ( .A(writeIn[83]), .Y(n579) );
  INVX2TS U914 ( .A(n579), .Y(n1714) );
  INVX2TS U915 ( .A(n579), .Y(n1715) );
  INVX2TS U916 ( .A(writeIn[84]), .Y(n580) );
  INVX2TS U917 ( .A(n580), .Y(n1716) );
  INVX2TS U918 ( .A(n580), .Y(n1717) );
  INVX2TS U919 ( .A(writeIn[85]), .Y(n581) );
  INVX2TS U920 ( .A(n581), .Y(n1718) );
  INVX2TS U921 ( .A(n581), .Y(n1719) );
  INVX2TS U922 ( .A(writeIn[86]), .Y(n582) );
  INVX2TS U923 ( .A(n582), .Y(n1720) );
  INVX2TS U924 ( .A(n582), .Y(n1721) );
  INVX2TS U925 ( .A(writeIn[87]), .Y(n583) );
  INVX2TS U926 ( .A(n583), .Y(n1722) );
  INVX2TS U927 ( .A(n583), .Y(n1723) );
  INVX2TS U928 ( .A(writeIn[88]), .Y(n584) );
  INVX2TS U929 ( .A(n584), .Y(n1724) );
  INVX2TS U930 ( .A(n584), .Y(n1725) );
  INVX2TS U931 ( .A(writeIn[89]), .Y(n585) );
  INVX2TS U932 ( .A(n585), .Y(n1726) );
  INVX2TS U933 ( .A(n585), .Y(n1727) );
  INVX2TS U934 ( .A(writeIn[90]), .Y(n586) );
  INVX2TS U935 ( .A(n586), .Y(n1728) );
  INVX2TS U936 ( .A(n586), .Y(n1729) );
  INVX2TS U937 ( .A(writeIn[91]), .Y(n587) );
  INVX2TS U938 ( .A(n587), .Y(n1730) );
  INVX2TS U939 ( .A(n587), .Y(n1731) );
  INVX2TS U940 ( .A(writeIn[92]), .Y(n588) );
  INVX2TS U941 ( .A(n588), .Y(n1732) );
  INVX2TS U942 ( .A(n588), .Y(n1733) );
  INVX2TS U943 ( .A(writeIn[93]), .Y(n589) );
  INVX2TS U944 ( .A(n589), .Y(n1734) );
  INVX2TS U945 ( .A(n589), .Y(n1735) );
  INVX2TS U946 ( .A(writeIn[94]), .Y(n590) );
  INVX2TS U947 ( .A(n590), .Y(n1736) );
  INVX2TS U948 ( .A(n590), .Y(n1737) );
  INVX2TS U949 ( .A(writeIn[95]), .Y(n591) );
  INVX2TS U950 ( .A(n591), .Y(n1738) );
  INVX2TS U951 ( .A(n591), .Y(n1739) );
  INVX2TS U952 ( .A(writeIn[96]), .Y(n592) );
  INVX2TS U953 ( .A(n592), .Y(n1740) );
  INVX2TS U954 ( .A(n592), .Y(n1741) );
  INVX2TS U955 ( .A(writeIn[97]), .Y(n593) );
  INVX2TS U956 ( .A(n593), .Y(n1742) );
  INVX2TS U957 ( .A(n593), .Y(n1743) );
  INVX2TS U958 ( .A(writeIn[98]), .Y(n594) );
  INVX2TS U959 ( .A(n594), .Y(n1744) );
  INVX2TS U960 ( .A(n594), .Y(n1745) );
  INVX2TS U961 ( .A(writeIn[99]), .Y(n595) );
  INVX2TS U962 ( .A(n595), .Y(n1746) );
  INVX2TS U963 ( .A(n595), .Y(n1747) );
  INVX2TS U964 ( .A(writeIn[100]), .Y(n596) );
  INVX2TS U965 ( .A(n596), .Y(n1748) );
  INVX2TS U966 ( .A(n596), .Y(n1749) );
  INVX2TS U967 ( .A(writeIn[101]), .Y(n597) );
  INVX2TS U968 ( .A(n597), .Y(n1750) );
  INVX2TS U969 ( .A(n597), .Y(n1751) );
  INVX2TS U970 ( .A(writeIn[102]), .Y(n598) );
  INVX2TS U971 ( .A(n598), .Y(n1752) );
  INVX2TS U972 ( .A(n598), .Y(n1753) );
  INVX2TS U973 ( .A(writeIn[103]), .Y(n599) );
  INVX2TS U974 ( .A(n599), .Y(n1754) );
  INVX2TS U975 ( .A(n599), .Y(n1755) );
  INVX2TS U976 ( .A(writeIn[104]), .Y(n600) );
  INVX2TS U977 ( .A(n600), .Y(n1756) );
  INVX2TS U978 ( .A(n600), .Y(n1757) );
  INVX2TS U979 ( .A(writeIn[105]), .Y(n601) );
  INVX2TS U980 ( .A(n601), .Y(n1758) );
  INVX2TS U981 ( .A(n601), .Y(n1759) );
  INVX2TS U982 ( .A(writeIn[106]), .Y(n602) );
  INVX2TS U983 ( .A(n602), .Y(n1760) );
  INVX2TS U984 ( .A(n602), .Y(n1761) );
  INVX2TS U985 ( .A(writeIn[107]), .Y(n603) );
  INVX2TS U986 ( .A(n603), .Y(n1762) );
  INVX2TS U987 ( .A(n603), .Y(n1763) );
  INVX2TS U988 ( .A(writeIn[108]), .Y(n604) );
  INVX2TS U989 ( .A(n604), .Y(n1764) );
  INVX2TS U990 ( .A(n604), .Y(n1765) );
  INVX2TS U991 ( .A(writeIn[109]), .Y(n605) );
  INVX2TS U992 ( .A(n605), .Y(n1766) );
  INVX2TS U993 ( .A(n605), .Y(n1767) );
  INVX2TS U994 ( .A(writeIn[110]), .Y(n606) );
  INVX2TS U995 ( .A(n606), .Y(n1768) );
  INVX2TS U996 ( .A(n606), .Y(n1769) );
  INVX2TS U997 ( .A(writeIn[111]), .Y(n607) );
  INVX2TS U998 ( .A(n607), .Y(n1770) );
  INVX2TS U999 ( .A(n607), .Y(n1771) );
  INVX2TS U1000 ( .A(writeIn[112]), .Y(n608) );
  INVX2TS U1001 ( .A(n608), .Y(n1772) );
  INVX2TS U1002 ( .A(n608), .Y(n1773) );
  INVX2TS U1003 ( .A(writeIn[113]), .Y(n609) );
  INVX2TS U1004 ( .A(n609), .Y(n1774) );
  INVX2TS U1005 ( .A(n609), .Y(n1775) );
  INVX2TS U1006 ( .A(writeIn[114]), .Y(n610) );
  INVX2TS U1007 ( .A(n610), .Y(n1776) );
  INVX2TS U1008 ( .A(n610), .Y(n1777) );
  INVX2TS U1009 ( .A(writeIn[115]), .Y(n611) );
  INVX2TS U1010 ( .A(n611), .Y(n1778) );
  INVX2TS U1011 ( .A(n611), .Y(n1779) );
  INVX2TS U1012 ( .A(writeIn[116]), .Y(n612) );
  INVX2TS U1013 ( .A(n612), .Y(n1780) );
  INVX2TS U1014 ( .A(n612), .Y(n1781) );
  INVX2TS U1015 ( .A(writeIn[117]), .Y(n613) );
  INVX2TS U1016 ( .A(n613), .Y(n1782) );
  INVX2TS U1017 ( .A(n613), .Y(n1783) );
  INVX2TS U1018 ( .A(writeIn[118]), .Y(n614) );
  INVX2TS U1019 ( .A(n614), .Y(n1784) );
  INVX2TS U1020 ( .A(n614), .Y(n1785) );
  INVX2TS U1021 ( .A(writeIn[119]), .Y(n615) );
  INVX2TS U1022 ( .A(n615), .Y(n1786) );
  INVX2TS U1023 ( .A(n615), .Y(n1787) );
  INVX2TS U1024 ( .A(writeIn[120]), .Y(n616) );
  INVX2TS U1025 ( .A(n616), .Y(n1788) );
  INVX2TS U1026 ( .A(n616), .Y(n1789) );
  INVX2TS U1027 ( .A(writeIn[121]), .Y(n617) );
  INVX2TS U1028 ( .A(n617), .Y(n1790) );
  INVX2TS U1029 ( .A(n617), .Y(n1791) );
  INVX2TS U1030 ( .A(writeIn[122]), .Y(n618) );
  INVX2TS U1031 ( .A(n618), .Y(n1792) );
  INVX2TS U1032 ( .A(n618), .Y(n1793) );
  INVX2TS U1033 ( .A(writeIn[123]), .Y(n619) );
  INVX2TS U1034 ( .A(n619), .Y(n1794) );
  INVX2TS U1035 ( .A(n619), .Y(n1795) );
  INVX2TS U1036 ( .A(writeIn[124]), .Y(n620) );
  INVX2TS U1037 ( .A(n620), .Y(n1796) );
  INVX2TS U1038 ( .A(n620), .Y(n1797) );
  INVX2TS U1039 ( .A(writeIn[125]), .Y(n621) );
  INVX2TS U1040 ( .A(n621), .Y(n1798) );
  INVX2TS U1041 ( .A(n621), .Y(n1799) );
  INVX2TS U1042 ( .A(writeIn[126]), .Y(n622) );
  INVX2TS U1043 ( .A(n622), .Y(n1800) );
  INVX2TS U1044 ( .A(n622), .Y(n1801) );
  INVX2TS U1045 ( .A(writeIn[127]), .Y(n623) );
  INVX2TS U1046 ( .A(n623), .Y(n1802) );
  INVX2TS U1047 ( .A(n623), .Y(n1803) );
  INVX2TS U1048 ( .A(writeIn[128]), .Y(n624) );
  INVX2TS U1049 ( .A(n624), .Y(n1804) );
  INVX2TS U1050 ( .A(n624), .Y(n1805) );
  INVX2TS U1051 ( .A(writeIn[129]), .Y(n625) );
  INVX2TS U1052 ( .A(n625), .Y(n1806) );
  INVX2TS U1053 ( .A(n625), .Y(n1807) );
  INVX2TS U1054 ( .A(writeIn[130]), .Y(n626) );
  INVX2TS U1055 ( .A(n626), .Y(n1808) );
  INVX2TS U1056 ( .A(n626), .Y(n1809) );
  INVX2TS U1057 ( .A(writeIn[131]), .Y(n627) );
  INVX2TS U1058 ( .A(n627), .Y(n1810) );
  INVX2TS U1059 ( .A(n627), .Y(n1811) );
  INVX2TS U1060 ( .A(writeIn[132]), .Y(n628) );
  INVX2TS U1061 ( .A(n628), .Y(n1812) );
  INVX2TS U1062 ( .A(n628), .Y(n1813) );
  INVX2TS U1063 ( .A(writeIn[133]), .Y(n629) );
  INVX2TS U1064 ( .A(n629), .Y(n1814) );
  INVX2TS U1065 ( .A(n629), .Y(n1815) );
  INVX2TS U1066 ( .A(writeIn[134]), .Y(n630) );
  INVX2TS U1067 ( .A(n630), .Y(n1816) );
  INVX2TS U1068 ( .A(n630), .Y(n1817) );
  INVX2TS U1069 ( .A(writeIn[135]), .Y(n631) );
  INVX2TS U1070 ( .A(n631), .Y(n1818) );
  INVX2TS U1071 ( .A(n631), .Y(n1819) );
  INVX2TS U1072 ( .A(writeIn[136]), .Y(n632) );
  INVX2TS U1073 ( .A(n632), .Y(n1820) );
  INVX2TS U1074 ( .A(n632), .Y(n1821) );
  INVX2TS U1075 ( .A(writeIn[137]), .Y(n633) );
  INVX2TS U1076 ( .A(n633), .Y(n1822) );
  INVX2TS U1077 ( .A(n633), .Y(n1823) );
  INVX2TS U1078 ( .A(writeIn[138]), .Y(n634) );
  INVX2TS U1079 ( .A(n634), .Y(n1824) );
  INVX2TS U1080 ( .A(n634), .Y(n1825) );
  INVX2TS U1081 ( .A(writeIn[139]), .Y(n635) );
  INVX2TS U1082 ( .A(n635), .Y(n1826) );
  INVX2TS U1083 ( .A(n635), .Y(n1827) );
  INVX2TS U1084 ( .A(writeIn[140]), .Y(n636) );
  INVX2TS U1085 ( .A(n636), .Y(n1828) );
  INVX2TS U1086 ( .A(n636), .Y(n1829) );
  INVX2TS U1087 ( .A(writeIn[141]), .Y(n637) );
  INVX2TS U1088 ( .A(n637), .Y(n1830) );
  INVX2TS U1089 ( .A(n637), .Y(n1831) );
  INVX2TS U1090 ( .A(writeIn[142]), .Y(n638) );
  INVX2TS U1091 ( .A(n638), .Y(n1832) );
  INVX2TS U1092 ( .A(n638), .Y(n1833) );
  INVX2TS U1093 ( .A(writeIn[143]), .Y(n639) );
  INVX2TS U1094 ( .A(n639), .Y(n1834) );
  INVX2TS U1095 ( .A(n639), .Y(n1835) );
  INVX2TS U1096 ( .A(writeIn[144]), .Y(n640) );
  INVX2TS U1097 ( .A(n640), .Y(n1836) );
  INVX2TS U1098 ( .A(n640), .Y(n1837) );
  INVX2TS U1099 ( .A(writeIn[145]), .Y(n641) );
  INVX2TS U1100 ( .A(n641), .Y(n1838) );
  INVX2TS U1101 ( .A(n641), .Y(n1839) );
  INVX2TS U1102 ( .A(writeIn[146]), .Y(n642) );
  INVX2TS U1103 ( .A(n642), .Y(n1840) );
  INVX2TS U1104 ( .A(n642), .Y(n1841) );
  INVX2TS U1105 ( .A(writeIn[147]), .Y(n643) );
  INVX2TS U1106 ( .A(n643), .Y(n1842) );
  INVX2TS U1107 ( .A(n643), .Y(n1843) );
  INVX2TS U1108 ( .A(writeIn[148]), .Y(n644) );
  INVX2TS U1109 ( .A(n644), .Y(n1844) );
  INVX2TS U1110 ( .A(n644), .Y(n1845) );
  INVX2TS U1111 ( .A(writeIn[149]), .Y(n645) );
  INVX2TS U1112 ( .A(n645), .Y(n1846) );
  INVX2TS U1113 ( .A(n645), .Y(n1847) );
  INVX2TS U1114 ( .A(writeIn[150]), .Y(n646) );
  INVX2TS U1115 ( .A(n646), .Y(n1848) );
  INVX2TS U1116 ( .A(n646), .Y(n1849) );
  INVX2TS U1117 ( .A(writeIn[151]), .Y(n647) );
  INVX2TS U1118 ( .A(n647), .Y(n1850) );
  INVX2TS U1119 ( .A(n647), .Y(n1851) );
  INVX2TS U1120 ( .A(writeIn[152]), .Y(n648) );
  INVX2TS U1121 ( .A(n648), .Y(n1852) );
  INVX2TS U1122 ( .A(n648), .Y(n1853) );
  INVX2TS U1123 ( .A(writeIn[153]), .Y(n649) );
  INVX2TS U1124 ( .A(n649), .Y(n1854) );
  INVX2TS U1125 ( .A(n649), .Y(n1855) );
  INVX2TS U1126 ( .A(writeIn[154]), .Y(n650) );
  INVX2TS U1127 ( .A(n650), .Y(n1856) );
  INVX2TS U1128 ( .A(n650), .Y(n1857) );
  INVX2TS U1129 ( .A(writeIn[155]), .Y(n651) );
  INVX2TS U1130 ( .A(n651), .Y(n1858) );
  INVX2TS U1131 ( .A(n651), .Y(n1859) );
  INVX2TS U1132 ( .A(writeIn[156]), .Y(n652) );
  INVX2TS U1133 ( .A(n652), .Y(n1860) );
  INVX2TS U1134 ( .A(n652), .Y(n1861) );
  INVX2TS U1135 ( .A(writeIn[157]), .Y(n653) );
  INVX2TS U1136 ( .A(n653), .Y(n1862) );
  INVX2TS U1137 ( .A(n653), .Y(n1863) );
  INVX2TS U1138 ( .A(writeIn[158]), .Y(n654) );
  INVX2TS U1139 ( .A(n654), .Y(n1864) );
  INVX2TS U1140 ( .A(n654), .Y(n1865) );
  INVX2TS U1141 ( .A(writeIn[159]), .Y(n655) );
  INVX2TS U1142 ( .A(n655), .Y(n1866) );
  INVX2TS U1143 ( .A(n655), .Y(n1867) );
  INVX2TS U1144 ( .A(NodeSelect[2]), .Y(n659) );
  INVX2TS U1145 ( .A(n659), .Y(n664) );
  INVX2TS U1146 ( .A(NodeSelect[0]), .Y(n656) );
  INVX2TS U1147 ( .A(n656), .Y(n677) );
  CLKINVX1TS U1148 ( .A(NodeSelect[1]), .Y(n678) );
  NOR3XLTS U1149 ( .A(n664), .B(n677), .C(n678), .Y(n1519) );
  CLKBUFX2TS U1150 ( .A(n1519), .Y(n1102) );
  CLKBUFX2TS U1151 ( .A(n1102), .Y(n1510) );
  CLKBUFX2TS U1152 ( .A(n1510), .Y(n1183) );
  CLKBUFX2TS U1153 ( .A(n1183), .Y(n1543) );
  CLKBUFX2TS U1154 ( .A(n1543), .Y(n1534) );
  NOR4XLTS U1155 ( .A(NodeSelect[5]), .B(NodeSelect[4]), .C(NodeSelect[9]), 
        .D(NodeSelect[8]), .Y(n657) );
  NAND3BXLTS U1156 ( .AN(NodeSelect[6]), .B(writeEnable), .C(n657), .Y(n660)
         );
  NOR3XLTS U1157 ( .A(NodeSelect[3]), .B(NodeSelect[7]), .C(n660), .Y(n679) );
  CLKAND2X2TS U1158 ( .A(n1534), .B(n679), .Y(n726) );
  CLKBUFX2TS U1159 ( .A(n726), .Y(n673) );
  CLKBUFX2TS U1160 ( .A(n673), .Y(n728) );
  CLKBUFX2TS U1161 ( .A(n728), .Y(n672) );
  CLKBUFX2TS U1162 ( .A(n672), .Y(n658) );
  CLKBUFX2TS U1163 ( .A(n658), .Y(n1984) );
  CLKBUFX2TS U1164 ( .A(n658), .Y(n1986) );
  CLKBUFX2TS U1165 ( .A(n658), .Y(n1987) );
  CLKBUFX2TS U1166 ( .A(n658), .Y(n1988) );
  CLKBUFX2TS U1167 ( .A(n673), .Y(n1872) );
  NOR3XLTS U1168 ( .A(n664), .B(n677), .C(NodeSelect[1]), .Y(n1517) );
  CLKBUFX2TS U1169 ( .A(n1517), .Y(n1101) );
  CLKBUFX2TS U1170 ( .A(n1101), .Y(n1508) );
  CLKBUFX2TS U1171 ( .A(n1508), .Y(n1181) );
  CLKBUFX2TS U1172 ( .A(n1181), .Y(n1541) );
  CLKBUFX2TS U1173 ( .A(n1541), .Y(n1532) );
  NOR3XLTS U1174 ( .A(NodeSelect[3]), .B(NodeSelect[7]), .C(n660), .Y(n680) );
  CLKAND2X2TS U1175 ( .A(n1532), .B(n680), .Y(n729) );
  CLKBUFX2TS U1176 ( .A(n729), .Y(n700) );
  CLKBUFX2TS U1177 ( .A(n700), .Y(n730) );
  CLKBUFX2TS U1178 ( .A(n730), .Y(n661) );
  CLKBUFX2TS U1179 ( .A(n661), .Y(n1890) );
  CLKBUFX2TS U1180 ( .A(n661), .Y(n1892) );
  CLKBUFX2TS U1181 ( .A(n661), .Y(n1893) );
  CLKBUFX2TS U1182 ( .A(n661), .Y(n1894) );
  CLKBUFX2TS U1183 ( .A(n728), .Y(n670) );
  CLKBUFX2TS U1184 ( .A(n670), .Y(n1979) );
  CLKBUFX2TS U1185 ( .A(n729), .Y(n675) );
  CLKBUFX2TS U1186 ( .A(n675), .Y(n731) );
  CLKBUFX2TS U1187 ( .A(n731), .Y(n662) );
  CLKBUFX2TS U1188 ( .A(n662), .Y(n1900) );
  CLKBUFX2TS U1189 ( .A(n662), .Y(n1901) );
  CLKBUFX2TS U1190 ( .A(n662), .Y(n1902) );
  CLKBUFX2TS U1191 ( .A(n662), .Y(n1903) );
  CLKBUFX2TS U1192 ( .A(n731), .Y(n674) );
  CLKBUFX2TS U1193 ( .A(n674), .Y(n663) );
  CLKBUFX2TS U1194 ( .A(n663), .Y(n1908) );
  CLKBUFX2TS U1195 ( .A(n663), .Y(n1910) );
  CLKBUFX2TS U1196 ( .A(n663), .Y(n1911) );
  CLKBUFX2TS U1197 ( .A(n663), .Y(n1912) );
  CLKBUFX2TS U1198 ( .A(n675), .Y(n1868) );
  NOR2XLTS U1199 ( .A(n677), .B(n659), .Y(n1080) );
  CLKBUFX2TS U1200 ( .A(n1080), .Y(n1506) );
  CLKBUFX2TS U1201 ( .A(n1506), .Y(n1179) );
  CLKBUFX2TS U1202 ( .A(n1179), .Y(n1539) );
  CLKBUFX2TS U1203 ( .A(n1539), .Y(n1530) );
  NAND2X1TS U1204 ( .A(n680), .B(n678), .Y(n681) );
  NOR2BX1TS U1205 ( .AN(n1530), .B(n681), .Y(n698) );
  CLKBUFX2TS U1206 ( .A(n698), .Y(n709) );
  CLKBUFX2TS U1207 ( .A(n709), .Y(n667) );
  CLKBUFX2TS U1208 ( .A(n667), .Y(n2035) );
  CLKBUFX2TS U1209 ( .A(n698), .Y(n708) );
  CLKBUFX2TS U1210 ( .A(n708), .Y(n665) );
  CLKBUFX2TS U1211 ( .A(n665), .Y(n2042) );
  CLKBUFX2TS U1212 ( .A(n665), .Y(n2044) );
  CLKBUFX2TS U1213 ( .A(n665), .Y(n2045) );
  CLKBUFX2TS U1214 ( .A(n665), .Y(n2046) );
  CLKBUFX2TS U1215 ( .A(n709), .Y(n671) );
  CLKBUFX2TS U1216 ( .A(n671), .Y(n725) );
  CLKBUFX2TS U1217 ( .A(n725), .Y(n666) );
  CLKBUFX2TS U1218 ( .A(n666), .Y(n2052) );
  CLKBUFX2TS U1219 ( .A(n666), .Y(n2053) );
  CLKBUFX2TS U1220 ( .A(n666), .Y(n2054) );
  CLKBUFX2TS U1221 ( .A(n666), .Y(n2055) );
  CLKBUFX2TS U1222 ( .A(n667), .Y(n2056) );
  CLKBUFX2TS U1223 ( .A(n667), .Y(n2057) );
  CLKBUFX2TS U1224 ( .A(n667), .Y(n2058) );
  CLKBUFX2TS U1225 ( .A(n725), .Y(n676) );
  CLKBUFX2TS U1226 ( .A(n676), .Y(n668) );
  CLKBUFX2TS U1227 ( .A(n668), .Y(n2060) );
  CLKBUFX2TS U1228 ( .A(n668), .Y(n2062) );
  CLKBUFX2TS U1229 ( .A(n668), .Y(n2063) );
  CLKBUFX2TS U1230 ( .A(n668), .Y(n2064) );
  CLKBUFX2TS U1231 ( .A(n671), .Y(n1876) );
  CLKBUFX2TS U1232 ( .A(n726), .Y(n699) );
  CLKBUFX2TS U1233 ( .A(n699), .Y(n727) );
  CLKBUFX2TS U1234 ( .A(n727), .Y(n669) );
  CLKBUFX2TS U1235 ( .A(n669), .Y(n1966) );
  CLKBUFX2TS U1236 ( .A(n669), .Y(n1968) );
  CLKBUFX2TS U1237 ( .A(n669), .Y(n1969) );
  CLKBUFX2TS U1238 ( .A(n669), .Y(n1970) );
  CLKBUFX2TS U1239 ( .A(n670), .Y(n1976) );
  CLKBUFX2TS U1240 ( .A(n670), .Y(n1977) );
  CLKBUFX2TS U1241 ( .A(n670), .Y(n1978) );
  CLKBUFX2TS U1242 ( .A(n671), .Y(n2051) );
  CLKBUFX2TS U1243 ( .A(n671), .Y(n2059) );
  CLKBUFX2TS U1244 ( .A(n727), .Y(n704) );
  CLKBUFX2TS U1245 ( .A(n704), .Y(n1963) );
  CLKBUFX2TS U1246 ( .A(n704), .Y(n1964) );
  CLKBUFX2TS U1247 ( .A(n672), .Y(n1971) );
  CLKBUFX2TS U1248 ( .A(n672), .Y(n1972) );
  CLKBUFX2TS U1249 ( .A(n672), .Y(n1973) );
  CLKBUFX2TS U1250 ( .A(n673), .Y(n1975) );
  CLKBUFX2TS U1251 ( .A(n673), .Y(n1983) );
  CLKBUFX2TS U1252 ( .A(n730), .Y(n706) );
  CLKBUFX2TS U1253 ( .A(n706), .Y(n1887) );
  CLKBUFX2TS U1254 ( .A(n706), .Y(n1888) );
  CLKBUFX2TS U1255 ( .A(n674), .Y(n1895) );
  CLKBUFX2TS U1256 ( .A(n674), .Y(n1896) );
  CLKBUFX2TS U1257 ( .A(n674), .Y(n1897) );
  CLKBUFX2TS U1258 ( .A(n675), .Y(n1899) );
  CLKBUFX2TS U1259 ( .A(n675), .Y(n1907) );
  CLKBUFX2TS U1260 ( .A(n1876), .Y(n1877) );
  CLKBUFX2TS U1261 ( .A(n1877), .Y(n2068) );
  CLKBUFX2TS U1262 ( .A(n1877), .Y(n2069) );
  CLKBUFX2TS U1263 ( .A(n1872), .Y(n1873) );
  CLKBUFX2TS U1264 ( .A(n1873), .Y(n1992) );
  CLKBUFX2TS U1265 ( .A(n1873), .Y(n1993) );
  CLKBUFX2TS U1266 ( .A(n1868), .Y(n1869) );
  CLKBUFX2TS U1267 ( .A(n1869), .Y(n1916) );
  CLKBUFX2TS U1268 ( .A(n1869), .Y(n1917) );
  CLKBUFX2TS U1269 ( .A(n708), .Y(n710) );
  CLKBUFX2TS U1270 ( .A(n710), .Y(n2039) );
  CLKBUFX2TS U1271 ( .A(n710), .Y(n2040) );
  CLKBUFX2TS U1272 ( .A(n676), .Y(n2047) );
  CLKBUFX2TS U1273 ( .A(n676), .Y(n2048) );
  CLKBUFX2TS U1274 ( .A(n676), .Y(n2049) );
  NOR3XLTS U1275 ( .A(n664), .B(n656), .C(n678), .Y(n1081) );
  CLKBUFX2TS U1276 ( .A(n1081), .Y(n818) );
  CLKBUFX2TS U1277 ( .A(n818), .Y(n1358) );
  CLKBUFX2TS U1278 ( .A(n1358), .Y(n1542) );
  CLKBUFX2TS U1279 ( .A(n1542), .Y(n1533) );
  CLKAND2X2TS U1280 ( .A(n1533), .B(n679), .Y(n741) );
  CLKBUFX2TS U1281 ( .A(n741), .Y(n687) );
  CLKBUFX2TS U1282 ( .A(n687), .Y(n1874) );
  CLKBUFX2TS U1283 ( .A(n1874), .Y(n1875) );
  CLKBUFX2TS U1284 ( .A(n1875), .Y(n2030) );
  CLKBUFX2TS U1285 ( .A(n1875), .Y(n2031) );
  NOR3XLTS U1286 ( .A(n664), .B(NodeSelect[1]), .C(n656), .Y(n1082) );
  CLKBUFX2TS U1287 ( .A(n1082), .Y(n820) );
  CLKBUFX2TS U1288 ( .A(n820), .Y(n1360) );
  CLKBUFX2TS U1289 ( .A(n1360), .Y(n1544) );
  CLKBUFX2TS U1290 ( .A(n1544), .Y(n1535) );
  CLKAND2X2TS U1291 ( .A(n1535), .B(n680), .Y(n737) );
  CLKBUFX2TS U1292 ( .A(n737), .Y(n688) );
  CLKBUFX2TS U1293 ( .A(n688), .Y(n1870) );
  CLKBUFX2TS U1294 ( .A(n1870), .Y(n1871) );
  CLKBUFX2TS U1295 ( .A(n1871), .Y(n1954) );
  CLKBUFX2TS U1296 ( .A(n1871), .Y(n1955) );
  NOR2XLTS U1297 ( .A(n659), .B(n656), .Y(n1507) );
  CLKBUFX2TS U1298 ( .A(n1507), .Y(n840) );
  CLKBUFX2TS U1299 ( .A(n840), .Y(n816) );
  CLKBUFX2TS U1300 ( .A(n816), .Y(n1298) );
  CLKBUFX2TS U1301 ( .A(n1298), .Y(n1056) );
  CLKBUFX2TS U1302 ( .A(n1056), .Y(n1540) );
  CLKBUFX2TS U1303 ( .A(n1540), .Y(n1531) );
  NOR2BX1TS U1304 ( .AN(n1531), .B(n681), .Y(n701) );
  CLKBUFX2TS U1305 ( .A(n701), .Y(n714) );
  CLKBUFX2TS U1306 ( .A(n714), .Y(n684) );
  CLKBUFX2TS U1307 ( .A(n684), .Y(n2073) );
  CLKBUFX2TS U1308 ( .A(n701), .Y(n715) );
  CLKBUFX2TS U1309 ( .A(n715), .Y(n682) );
  CLKBUFX2TS U1310 ( .A(n682), .Y(n2080) );
  CLKBUFX2TS U1311 ( .A(n682), .Y(n2082) );
  CLKBUFX2TS U1312 ( .A(n682), .Y(n2083) );
  CLKBUFX2TS U1313 ( .A(n682), .Y(n2084) );
  CLKBUFX2TS U1314 ( .A(n714), .Y(n686) );
  CLKBUFX2TS U1315 ( .A(n686), .Y(n740) );
  CLKBUFX2TS U1316 ( .A(n740), .Y(n683) );
  CLKBUFX2TS U1317 ( .A(n683), .Y(n2090) );
  CLKBUFX2TS U1318 ( .A(n683), .Y(n2091) );
  CLKBUFX2TS U1319 ( .A(n683), .Y(n2092) );
  CLKBUFX2TS U1320 ( .A(n683), .Y(n2093) );
  CLKBUFX2TS U1321 ( .A(n684), .Y(n2094) );
  CLKBUFX2TS U1322 ( .A(n684), .Y(n2095) );
  CLKBUFX2TS U1323 ( .A(n684), .Y(n2096) );
  CLKBUFX2TS U1324 ( .A(n740), .Y(n693) );
  CLKBUFX2TS U1325 ( .A(n693), .Y(n685) );
  CLKBUFX2TS U1326 ( .A(n685), .Y(n2098) );
  CLKBUFX2TS U1327 ( .A(n685), .Y(n2100) );
  CLKBUFX2TS U1328 ( .A(n685), .Y(n2101) );
  CLKBUFX2TS U1329 ( .A(n685), .Y(n2102) );
  CLKBUFX2TS U1330 ( .A(n686), .Y(n1878) );
  CLKBUFX2TS U1331 ( .A(n1878), .Y(n1879) );
  CLKBUFX2TS U1332 ( .A(n1879), .Y(n2106) );
  CLKBUFX2TS U1333 ( .A(n1879), .Y(n2107) );
  CLKBUFX2TS U1334 ( .A(n693), .Y(n2087) );
  CLKBUFX2TS U1335 ( .A(n686), .Y(n2089) );
  CLKBUFX2TS U1336 ( .A(n686), .Y(n2097) );
  CLKBUFX2TS U1337 ( .A(n741), .Y(n702) );
  CLKBUFX2TS U1338 ( .A(n702), .Y(n742) );
  CLKBUFX2TS U1339 ( .A(n742), .Y(n716) );
  CLKBUFX2TS U1340 ( .A(n716), .Y(n2001) );
  CLKBUFX2TS U1341 ( .A(n716), .Y(n2002) );
  CLKBUFX2TS U1342 ( .A(n687), .Y(n743) );
  CLKBUFX2TS U1343 ( .A(n743), .Y(n691) );
  CLKBUFX2TS U1344 ( .A(n691), .Y(n2009) );
  CLKBUFX2TS U1345 ( .A(n691), .Y(n2010) );
  CLKBUFX2TS U1346 ( .A(n691), .Y(n2011) );
  CLKBUFX2TS U1347 ( .A(n687), .Y(n2013) );
  CLKBUFX2TS U1348 ( .A(n687), .Y(n2021) );
  CLKBUFX2TS U1349 ( .A(n737), .Y(n703) );
  CLKBUFX2TS U1350 ( .A(n703), .Y(n732) );
  CLKBUFX2TS U1351 ( .A(n732), .Y(n717) );
  CLKBUFX2TS U1352 ( .A(n717), .Y(n1925) );
  CLKBUFX2TS U1353 ( .A(n717), .Y(n1926) );
  CLKBUFX2TS U1354 ( .A(n688), .Y(n733) );
  CLKBUFX2TS U1355 ( .A(n733), .Y(n694) );
  CLKBUFX2TS U1356 ( .A(n694), .Y(n1933) );
  CLKBUFX2TS U1357 ( .A(n694), .Y(n1934) );
  CLKBUFX2TS U1358 ( .A(n694), .Y(n1935) );
  CLKBUFX2TS U1359 ( .A(n688), .Y(n1937) );
  CLKBUFX2TS U1360 ( .A(n688), .Y(n1945) );
  CLKBUFX2TS U1361 ( .A(n742), .Y(n689) );
  CLKBUFX2TS U1362 ( .A(n689), .Y(n2004) );
  CLKBUFX2TS U1363 ( .A(n689), .Y(n2006) );
  CLKBUFX2TS U1364 ( .A(n689), .Y(n2007) );
  CLKBUFX2TS U1365 ( .A(n689), .Y(n2008) );
  CLKBUFX2TS U1366 ( .A(n743), .Y(n690) );
  CLKBUFX2TS U1367 ( .A(n690), .Y(n2014) );
  CLKBUFX2TS U1368 ( .A(n690), .Y(n2015) );
  CLKBUFX2TS U1369 ( .A(n690), .Y(n2016) );
  CLKBUFX2TS U1370 ( .A(n690), .Y(n2017) );
  CLKBUFX2TS U1371 ( .A(n691), .Y(n692) );
  CLKBUFX2TS U1372 ( .A(n692), .Y(n2022) );
  CLKBUFX2TS U1373 ( .A(n692), .Y(n2024) );
  CLKBUFX2TS U1374 ( .A(n692), .Y(n2025) );
  CLKBUFX2TS U1375 ( .A(n692), .Y(n2026) );
  CLKBUFX2TS U1376 ( .A(n732), .Y(n697) );
  CLKBUFX2TS U1377 ( .A(n697), .Y(n1928) );
  CLKBUFX2TS U1378 ( .A(n693), .Y(n2086) );
  CLKBUFX2TS U1379 ( .A(n693), .Y(n2085) );
  CLKBUFX2TS U1380 ( .A(n715), .Y(n712) );
  CLKBUFX2TS U1381 ( .A(n712), .Y(n2078) );
  CLKBUFX2TS U1382 ( .A(n712), .Y(n2077) );
  CLKBUFX2TS U1383 ( .A(n694), .Y(n695) );
  CLKBUFX2TS U1384 ( .A(n695), .Y(n1950) );
  CLKBUFX2TS U1385 ( .A(n695), .Y(n1949) );
  CLKBUFX2TS U1386 ( .A(n695), .Y(n1948) );
  CLKBUFX2TS U1387 ( .A(n695), .Y(n1946) );
  CLKBUFX2TS U1388 ( .A(n733), .Y(n696) );
  CLKBUFX2TS U1389 ( .A(n696), .Y(n1941) );
  CLKBUFX2TS U1390 ( .A(n696), .Y(n1940) );
  CLKBUFX2TS U1391 ( .A(n696), .Y(n1939) );
  CLKBUFX2TS U1392 ( .A(n696), .Y(n1938) );
  CLKBUFX2TS U1393 ( .A(n697), .Y(n1932) );
  CLKBUFX2TS U1394 ( .A(n697), .Y(n1931) );
  CLKBUFX2TS U1395 ( .A(n697), .Y(n1930) );
  CLKBUFX2TS U1396 ( .A(n698), .Y(n2038) );
  CLKBUFX2TS U1397 ( .A(n699), .Y(n1957) );
  CLKBUFX2TS U1398 ( .A(n699), .Y(n1959) );
  CLKBUFX2TS U1399 ( .A(n699), .Y(n1962) );
  CLKBUFX2TS U1400 ( .A(n700), .Y(n1881) );
  CLKBUFX2TS U1401 ( .A(n700), .Y(n1883) );
  CLKBUFX2TS U1402 ( .A(n700), .Y(n1886) );
  CLKBUFX2TS U1403 ( .A(n701), .Y(n2076) );
  CLKBUFX2TS U1404 ( .A(n702), .Y(n1995) );
  CLKBUFX2TS U1405 ( .A(n702), .Y(n1997) );
  CLKBUFX2TS U1406 ( .A(n702), .Y(n2000) );
  CLKBUFX2TS U1407 ( .A(n703), .Y(n1919) );
  CLKBUFX2TS U1408 ( .A(n703), .Y(n1921) );
  CLKBUFX2TS U1409 ( .A(n703), .Y(n1924) );
  CLKBUFX2TS U1410 ( .A(n709), .Y(n2033) );
  CLKBUFX2TS U1411 ( .A(n704), .Y(n705) );
  CLKBUFX2TS U1412 ( .A(n705), .Y(n1956) );
  CLKBUFX2TS U1413 ( .A(n705), .Y(n1960) );
  CLKBUFX2TS U1414 ( .A(n705), .Y(n1961) );
  CLKBUFX2TS U1415 ( .A(n706), .Y(n707) );
  CLKBUFX2TS U1416 ( .A(n707), .Y(n1880) );
  CLKBUFX2TS U1417 ( .A(n707), .Y(n1884) );
  CLKBUFX2TS U1418 ( .A(n707), .Y(n1885) );
  CLKBUFX2TS U1419 ( .A(n708), .Y(n2041) );
  CLKBUFX2TS U1420 ( .A(n708), .Y(n2043) );
  CLKBUFX2TS U1421 ( .A(n709), .Y(n2034) );
  CLKBUFX2TS U1422 ( .A(n710), .Y(n711) );
  CLKBUFX2TS U1423 ( .A(n711), .Y(n2032) );
  CLKBUFX2TS U1424 ( .A(n711), .Y(n2036) );
  CLKBUFX2TS U1425 ( .A(n711), .Y(n2037) );
  CLKBUFX2TS U1426 ( .A(n712), .Y(n713) );
  CLKBUFX2TS U1427 ( .A(n713), .Y(n2070) );
  CLKBUFX2TS U1428 ( .A(n713), .Y(n2074) );
  CLKBUFX2TS U1429 ( .A(n713), .Y(n2075) );
  CLKBUFX2TS U1430 ( .A(n714), .Y(n2071) );
  CLKBUFX2TS U1431 ( .A(n714), .Y(n2072) );
  CLKBUFX2TS U1432 ( .A(n715), .Y(n2079) );
  CLKBUFX2TS U1433 ( .A(n715), .Y(n2081) );
  CLKBUFX2TS U1434 ( .A(n716), .Y(n718) );
  CLKBUFX2TS U1435 ( .A(n718), .Y(n1998) );
  CLKBUFX2TS U1436 ( .A(n718), .Y(n1999) );
  CLKBUFX2TS U1437 ( .A(n717), .Y(n719) );
  CLKBUFX2TS U1438 ( .A(n719), .Y(n1922) );
  CLKBUFX2TS U1439 ( .A(n719), .Y(n1923) );
  CLKBUFX2TS U1440 ( .A(n718), .Y(n1994) );
  CLKBUFX2TS U1441 ( .A(n719), .Y(n1918) );
  CLKBUFX2TS U1442 ( .A(n726), .Y(n720) );
  CLKBUFX2TS U1443 ( .A(n720), .Y(n1980) );
  CLKBUFX2TS U1444 ( .A(n720), .Y(n1981) );
  CLKBUFX2TS U1445 ( .A(n720), .Y(n1982) );
  CLKBUFX2TS U1446 ( .A(n1872), .Y(n721) );
  CLKBUFX2TS U1447 ( .A(n721), .Y(n1989) );
  CLKBUFX2TS U1448 ( .A(n721), .Y(n1990) );
  CLKBUFX2TS U1449 ( .A(n721), .Y(n1991) );
  CLKBUFX2TS U1450 ( .A(n729), .Y(n722) );
  CLKBUFX2TS U1451 ( .A(n722), .Y(n1904) );
  CLKBUFX2TS U1452 ( .A(n722), .Y(n1905) );
  CLKBUFX2TS U1453 ( .A(n722), .Y(n1906) );
  CLKBUFX2TS U1454 ( .A(n1868), .Y(n723) );
  CLKBUFX2TS U1455 ( .A(n723), .Y(n1913) );
  CLKBUFX2TS U1456 ( .A(n723), .Y(n1914) );
  CLKBUFX2TS U1457 ( .A(n723), .Y(n1915) );
  CLKBUFX2TS U1458 ( .A(n1876), .Y(n724) );
  CLKBUFX2TS U1459 ( .A(n724), .Y(n2065) );
  CLKBUFX2TS U1460 ( .A(n724), .Y(n2066) );
  CLKBUFX2TS U1461 ( .A(n724), .Y(n2067) );
  CLKBUFX2TS U1462 ( .A(n725), .Y(n2050) );
  CLKBUFX2TS U1463 ( .A(n725), .Y(n2061) );
  CLKBUFX2TS U1464 ( .A(n726), .Y(n1958) );
  CLKBUFX2TS U1465 ( .A(n727), .Y(n1965) );
  CLKBUFX2TS U1466 ( .A(n727), .Y(n1967) );
  CLKBUFX2TS U1467 ( .A(n728), .Y(n1974) );
  CLKBUFX2TS U1468 ( .A(n728), .Y(n1985) );
  CLKBUFX2TS U1469 ( .A(n729), .Y(n1882) );
  CLKBUFX2TS U1470 ( .A(n730), .Y(n1889) );
  CLKBUFX2TS U1471 ( .A(n730), .Y(n1891) );
  CLKBUFX2TS U1472 ( .A(n731), .Y(n1898) );
  CLKBUFX2TS U1473 ( .A(n731), .Y(n1909) );
  CLKBUFX2TS U1474 ( .A(n743), .Y(n2023) );
  CLKBUFX2TS U1475 ( .A(n737), .Y(n1920) );
  CLKBUFX2TS U1476 ( .A(n732), .Y(n1927) );
  CLKBUFX2TS U1477 ( .A(n732), .Y(n1929) );
  CLKBUFX2TS U1478 ( .A(n733), .Y(n1936) );
  CLKBUFX2TS U1479 ( .A(n733), .Y(n1947) );
  CLKBUFX2TS U1480 ( .A(n1878), .Y(n734) );
  CLKBUFX2TS U1481 ( .A(n734), .Y(n2103) );
  CLKBUFX2TS U1482 ( .A(n734), .Y(n2104) );
  CLKBUFX2TS U1483 ( .A(n734), .Y(n2105) );
  CLKBUFX2TS U1484 ( .A(n741), .Y(n735) );
  CLKBUFX2TS U1485 ( .A(n735), .Y(n2018) );
  CLKBUFX2TS U1486 ( .A(n735), .Y(n2019) );
  CLKBUFX2TS U1487 ( .A(n735), .Y(n2020) );
  CLKBUFX2TS U1488 ( .A(n1874), .Y(n736) );
  CLKBUFX2TS U1489 ( .A(n736), .Y(n2027) );
  CLKBUFX2TS U1490 ( .A(n736), .Y(n2028) );
  CLKBUFX2TS U1491 ( .A(n736), .Y(n2029) );
  CLKBUFX2TS U1492 ( .A(n737), .Y(n738) );
  CLKBUFX2TS U1493 ( .A(n738), .Y(n1942) );
  CLKBUFX2TS U1494 ( .A(n738), .Y(n1943) );
  CLKBUFX2TS U1495 ( .A(n738), .Y(n1944) );
  CLKBUFX2TS U1496 ( .A(n1870), .Y(n739) );
  CLKBUFX2TS U1497 ( .A(n739), .Y(n1951) );
  CLKBUFX2TS U1498 ( .A(n739), .Y(n1952) );
  CLKBUFX2TS U1499 ( .A(n739), .Y(n1953) );
  CLKBUFX2TS U1500 ( .A(n740), .Y(n2088) );
  CLKBUFX2TS U1501 ( .A(n740), .Y(n2099) );
  CLKBUFX2TS U1502 ( .A(n741), .Y(n1996) );
  CLKBUFX2TS U1503 ( .A(n742), .Y(n2003) );
  CLKBUFX2TS U1504 ( .A(n742), .Y(n2005) );
  CLKBUFX2TS U1505 ( .A(n743), .Y(n2012) );
  CLKBUFX2TS U1506 ( .A(n840), .Y(n756) );
  CLKBUFX2TS U1507 ( .A(n1506), .Y(n1299) );
  CLKBUFX2TS U1508 ( .A(n1299), .Y(n1477) );
  CLKBUFX2TS U1509 ( .A(n1477), .Y(n1239) );
  CLKBUFX2TS U1510 ( .A(n1239), .Y(n841) );
  CLKBUFX2TS U1511 ( .A(n841), .Y(n757) );
  AOI22X1TS U1512 ( .A0(n756), .A1(readOutBus[959]), .B0(n757), .B1(
        readOutBus[799]), .Y(n746) );
  CLKBUFX2TS U1513 ( .A(n1081), .Y(n1509) );
  CLKBUFX2TS U1514 ( .A(n1509), .Y(n758) );
  CLKBUFX2TS U1515 ( .A(n1508), .Y(n1300) );
  CLKBUFX2TS U1516 ( .A(n1300), .Y(n1479) );
  CLKBUFX2TS U1517 ( .A(n1479), .Y(n1241) );
  CLKBUFX2TS U1518 ( .A(n1241), .Y(n842) );
  CLKBUFX2TS U1519 ( .A(n842), .Y(n759) );
  AOI22X1TS U1520 ( .A0(n758), .A1(readOutBus[639]), .B0(n759), .B1(
        readOutBus[159]), .Y(n745) );
  CLKBUFX2TS U1521 ( .A(n1082), .Y(n1511) );
  CLKBUFX2TS U1522 ( .A(n1511), .Y(n760) );
  CLKBUFX2TS U1523 ( .A(n1510), .Y(n1301) );
  CLKBUFX2TS U1524 ( .A(n1301), .Y(n1481) );
  CLKBUFX2TS U1525 ( .A(n1481), .Y(n1243) );
  CLKBUFX2TS U1526 ( .A(n1243), .Y(n843) );
  CLKBUFX2TS U1527 ( .A(n843), .Y(n761) );
  AOI22X1TS U1528 ( .A0(n760), .A1(readOutBus[319]), .B0(n761), .B1(
        readOutBus[479]), .Y(n744) );
  NAND3XLTS U1529 ( .A(n746), .B(n745), .C(n744), .Y(readOut[159]) );
  AOI22X1TS U1530 ( .A0(n756), .A1(readOutBus[958]), .B0(n757), .B1(
        readOutBus[798]), .Y(n749) );
  AOI22X1TS U1531 ( .A0(n758), .A1(readOutBus[638]), .B0(n759), .B1(
        readOutBus[158]), .Y(n748) );
  AOI22X1TS U1532 ( .A0(n760), .A1(readOutBus[318]), .B0(n761), .B1(
        readOutBus[478]), .Y(n747) );
  NAND3XLTS U1533 ( .A(n749), .B(n748), .C(n747), .Y(readOut[158]) );
  AOI22X1TS U1534 ( .A0(n756), .A1(readOutBus[957]), .B0(n757), .B1(
        readOutBus[797]), .Y(n752) );
  AOI22X1TS U1535 ( .A0(n758), .A1(readOutBus[637]), .B0(n759), .B1(
        readOutBus[157]), .Y(n751) );
  AOI22X1TS U1536 ( .A0(n760), .A1(readOutBus[317]), .B0(n761), .B1(
        readOutBus[477]), .Y(n750) );
  NAND3XLTS U1537 ( .A(n752), .B(n751), .C(n750), .Y(readOut[157]) );
  AOI22X1TS U1538 ( .A0(n840), .A1(readOutBus[956]), .B0(n841), .B1(
        readOutBus[796]), .Y(n755) );
  AOI22X1TS U1539 ( .A0(n1081), .A1(readOutBus[636]), .B0(n842), .B1(
        readOutBus[156]), .Y(n754) );
  AOI22X1TS U1540 ( .A0(n1082), .A1(readOutBus[316]), .B0(n843), .B1(
        readOutBus[476]), .Y(n753) );
  NAND3XLTS U1541 ( .A(n755), .B(n754), .C(n753), .Y(readOut[156]) );
  CLKBUFX2TS U1542 ( .A(n756), .Y(n772) );
  CLKBUFX2TS U1543 ( .A(n757), .Y(n771) );
  AOI22X1TS U1544 ( .A0(n772), .A1(readOutBus[955]), .B0(n771), .B1(
        readOutBus[795]), .Y(n764) );
  CLKBUFX2TS U1545 ( .A(n758), .Y(n774) );
  CLKBUFX2TS U1546 ( .A(n759), .Y(n773) );
  AOI22X1TS U1547 ( .A0(n774), .A1(readOutBus[635]), .B0(n773), .B1(
        readOutBus[155]), .Y(n763) );
  CLKBUFX2TS U1548 ( .A(n760), .Y(n776) );
  CLKBUFX2TS U1549 ( .A(n761), .Y(n775) );
  AOI22X1TS U1550 ( .A0(n776), .A1(readOutBus[315]), .B0(n775), .B1(
        readOutBus[475]), .Y(n762) );
  NAND3XLTS U1551 ( .A(n764), .B(n763), .C(n762), .Y(readOut[155]) );
  AOI22X1TS U1552 ( .A0(n772), .A1(readOutBus[954]), .B0(n771), .B1(
        readOutBus[794]), .Y(n767) );
  AOI22X1TS U1553 ( .A0(n774), .A1(readOutBus[634]), .B0(n773), .B1(
        readOutBus[154]), .Y(n766) );
  AOI22X1TS U1554 ( .A0(n776), .A1(readOutBus[314]), .B0(n775), .B1(
        readOutBus[474]), .Y(n765) );
  NAND3XLTS U1555 ( .A(n767), .B(n766), .C(n765), .Y(readOut[154]) );
  AOI22X1TS U1556 ( .A0(n772), .A1(readOutBus[953]), .B0(n771), .B1(
        readOutBus[793]), .Y(n770) );
  AOI22X1TS U1557 ( .A0(n774), .A1(readOutBus[633]), .B0(n773), .B1(
        readOutBus[153]), .Y(n769) );
  AOI22X1TS U1558 ( .A0(n776), .A1(readOutBus[313]), .B0(n775), .B1(
        readOutBus[473]), .Y(n768) );
  NAND3XLTS U1559 ( .A(n770), .B(n769), .C(n768), .Y(readOut[153]) );
  AOI22X1TS U1560 ( .A0(n772), .A1(readOutBus[952]), .B0(n771), .B1(
        readOutBus[792]), .Y(n779) );
  AOI22X1TS U1561 ( .A0(n774), .A1(readOutBus[632]), .B0(n773), .B1(
        readOutBus[152]), .Y(n778) );
  AOI22X1TS U1562 ( .A0(n776), .A1(readOutBus[312]), .B0(n775), .B1(
        readOutBus[472]), .Y(n777) );
  NAND3XLTS U1563 ( .A(n779), .B(n778), .C(n777), .Y(readOut[152]) );
  CLKBUFX2TS U1564 ( .A(n816), .Y(n790) );
  CLKBUFX2TS U1565 ( .A(n841), .Y(n817) );
  CLKBUFX2TS U1566 ( .A(n817), .Y(n789) );
  AOI22X1TS U1567 ( .A0(n790), .A1(readOutBus[951]), .B0(n789), .B1(
        readOutBus[791]), .Y(n782) );
  CLKBUFX2TS U1568 ( .A(n818), .Y(n792) );
  CLKBUFX2TS U1569 ( .A(n842), .Y(n819) );
  CLKBUFX2TS U1570 ( .A(n819), .Y(n791) );
  AOI22X1TS U1571 ( .A0(n792), .A1(readOutBus[631]), .B0(n791), .B1(
        readOutBus[151]), .Y(n781) );
  CLKBUFX2TS U1572 ( .A(n820), .Y(n794) );
  CLKBUFX2TS U1573 ( .A(n843), .Y(n821) );
  CLKBUFX2TS U1574 ( .A(n821), .Y(n793) );
  AOI22X1TS U1575 ( .A0(n794), .A1(readOutBus[311]), .B0(n793), .B1(
        readOutBus[471]), .Y(n780) );
  NAND3XLTS U1576 ( .A(n782), .B(n781), .C(n780), .Y(readOut[151]) );
  AOI22X1TS U1577 ( .A0(n790), .A1(readOutBus[950]), .B0(n789), .B1(
        readOutBus[790]), .Y(n785) );
  AOI22X1TS U1578 ( .A0(n792), .A1(readOutBus[630]), .B0(n791), .B1(
        readOutBus[150]), .Y(n784) );
  AOI22X1TS U1579 ( .A0(n794), .A1(readOutBus[310]), .B0(n793), .B1(
        readOutBus[470]), .Y(n783) );
  NAND3XLTS U1580 ( .A(n785), .B(n784), .C(n783), .Y(readOut[150]) );
  AOI22X1TS U1581 ( .A0(n790), .A1(readOutBus[949]), .B0(n789), .B1(
        readOutBus[789]), .Y(n788) );
  AOI22X1TS U1582 ( .A0(n792), .A1(readOutBus[629]), .B0(n791), .B1(
        readOutBus[149]), .Y(n787) );
  AOI22X1TS U1583 ( .A0(n794), .A1(readOutBus[309]), .B0(n793), .B1(
        readOutBus[469]), .Y(n786) );
  NAND3XLTS U1584 ( .A(n788), .B(n787), .C(n786), .Y(readOut[149]) );
  AOI22X1TS U1585 ( .A0(n790), .A1(readOutBus[948]), .B0(n789), .B1(
        readOutBus[788]), .Y(n797) );
  AOI22X1TS U1586 ( .A0(n792), .A1(readOutBus[628]), .B0(n791), .B1(
        readOutBus[148]), .Y(n796) );
  AOI22X1TS U1587 ( .A0(n794), .A1(readOutBus[308]), .B0(n793), .B1(
        readOutBus[468]), .Y(n795) );
  NAND3XLTS U1588 ( .A(n797), .B(n796), .C(n795), .Y(readOut[148]) );
  CLKBUFX2TS U1589 ( .A(n816), .Y(n808) );
  CLKBUFX2TS U1590 ( .A(n817), .Y(n807) );
  AOI22X1TS U1591 ( .A0(n808), .A1(readOutBus[947]), .B0(n807), .B1(
        readOutBus[787]), .Y(n800) );
  CLKBUFX2TS U1592 ( .A(n818), .Y(n810) );
  CLKBUFX2TS U1593 ( .A(n819), .Y(n809) );
  AOI22X1TS U1594 ( .A0(n810), .A1(readOutBus[627]), .B0(n809), .B1(
        readOutBus[147]), .Y(n799) );
  CLKBUFX2TS U1595 ( .A(n820), .Y(n812) );
  CLKBUFX2TS U1596 ( .A(n821), .Y(n811) );
  AOI22X1TS U1597 ( .A0(n812), .A1(readOutBus[307]), .B0(n811), .B1(
        readOutBus[467]), .Y(n798) );
  NAND3XLTS U1598 ( .A(n800), .B(n799), .C(n798), .Y(readOut[147]) );
  AOI22X1TS U1599 ( .A0(n808), .A1(readOutBus[946]), .B0(n807), .B1(
        readOutBus[786]), .Y(n803) );
  AOI22X1TS U1600 ( .A0(n810), .A1(readOutBus[626]), .B0(n809), .B1(
        readOutBus[146]), .Y(n802) );
  AOI22X1TS U1601 ( .A0(n812), .A1(readOutBus[306]), .B0(n811), .B1(
        readOutBus[466]), .Y(n801) );
  NAND3XLTS U1602 ( .A(n803), .B(n802), .C(n801), .Y(readOut[146]) );
  AOI22X1TS U1603 ( .A0(n808), .A1(readOutBus[945]), .B0(n807), .B1(
        readOutBus[785]), .Y(n806) );
  AOI22X1TS U1604 ( .A0(n810), .A1(readOutBus[625]), .B0(n809), .B1(
        readOutBus[145]), .Y(n805) );
  AOI22X1TS U1605 ( .A0(n812), .A1(readOutBus[305]), .B0(n811), .B1(
        readOutBus[465]), .Y(n804) );
  NAND3XLTS U1606 ( .A(n806), .B(n805), .C(n804), .Y(readOut[145]) );
  AOI22X1TS U1607 ( .A0(n808), .A1(readOutBus[944]), .B0(n807), .B1(
        readOutBus[784]), .Y(n815) );
  AOI22X1TS U1608 ( .A0(n810), .A1(readOutBus[624]), .B0(n809), .B1(
        readOutBus[144]), .Y(n814) );
  AOI22X1TS U1609 ( .A0(n812), .A1(readOutBus[304]), .B0(n811), .B1(
        readOutBus[464]), .Y(n813) );
  NAND3XLTS U1610 ( .A(n815), .B(n814), .C(n813), .Y(readOut[144]) );
  CLKBUFX2TS U1611 ( .A(n816), .Y(n832) );
  CLKBUFX2TS U1612 ( .A(n817), .Y(n831) );
  AOI22X1TS U1613 ( .A0(n832), .A1(readOutBus[943]), .B0(n831), .B1(
        readOutBus[783]), .Y(n824) );
  CLKBUFX2TS U1614 ( .A(n818), .Y(n834) );
  CLKBUFX2TS U1615 ( .A(n819), .Y(n833) );
  AOI22X1TS U1616 ( .A0(n834), .A1(readOutBus[623]), .B0(n833), .B1(
        readOutBus[143]), .Y(n823) );
  CLKBUFX2TS U1617 ( .A(n820), .Y(n836) );
  CLKBUFX2TS U1618 ( .A(n821), .Y(n835) );
  AOI22X1TS U1619 ( .A0(n836), .A1(readOutBus[303]), .B0(n835), .B1(
        readOutBus[463]), .Y(n822) );
  NAND3XLTS U1620 ( .A(n824), .B(n823), .C(n822), .Y(readOut[143]) );
  AOI22X1TS U1621 ( .A0(n832), .A1(readOutBus[942]), .B0(n831), .B1(
        readOutBus[782]), .Y(n827) );
  AOI22X1TS U1622 ( .A0(n834), .A1(readOutBus[622]), .B0(n833), .B1(
        readOutBus[142]), .Y(n826) );
  AOI22X1TS U1623 ( .A0(n836), .A1(readOutBus[302]), .B0(n835), .B1(
        readOutBus[462]), .Y(n825) );
  NAND3XLTS U1624 ( .A(n827), .B(n826), .C(n825), .Y(readOut[142]) );
  AOI22X1TS U1625 ( .A0(n832), .A1(readOutBus[941]), .B0(n831), .B1(
        readOutBus[781]), .Y(n830) );
  AOI22X1TS U1626 ( .A0(n834), .A1(readOutBus[621]), .B0(n833), .B1(
        readOutBus[141]), .Y(n829) );
  AOI22X1TS U1627 ( .A0(n836), .A1(readOutBus[301]), .B0(n835), .B1(
        readOutBus[461]), .Y(n828) );
  NAND3XLTS U1628 ( .A(n830), .B(n829), .C(n828), .Y(readOut[141]) );
  AOI22X1TS U1629 ( .A0(n832), .A1(readOutBus[940]), .B0(n831), .B1(
        readOutBus[780]), .Y(n839) );
  AOI22X1TS U1630 ( .A0(n834), .A1(readOutBus[620]), .B0(n833), .B1(
        readOutBus[140]), .Y(n838) );
  AOI22X1TS U1631 ( .A0(n836), .A1(readOutBus[300]), .B0(n835), .B1(
        readOutBus[460]), .Y(n837) );
  NAND3XLTS U1632 ( .A(n839), .B(n838), .C(n837), .Y(readOut[140]) );
  CLKBUFX2TS U1633 ( .A(n840), .Y(n880) );
  CLKBUFX2TS U1634 ( .A(n880), .Y(n854) );
  CLKBUFX2TS U1635 ( .A(n841), .Y(n881) );
  CLKBUFX2TS U1636 ( .A(n881), .Y(n853) );
  AOI22X1TS U1637 ( .A0(n854), .A1(readOutBus[939]), .B0(n853), .B1(
        readOutBus[779]), .Y(n846) );
  CLKBUFX2TS U1638 ( .A(n1509), .Y(n902) );
  CLKBUFX2TS U1639 ( .A(n902), .Y(n856) );
  CLKBUFX2TS U1640 ( .A(n842), .Y(n882) );
  CLKBUFX2TS U1641 ( .A(n882), .Y(n855) );
  AOI22X1TS U1642 ( .A0(n856), .A1(readOutBus[619]), .B0(n855), .B1(
        readOutBus[139]), .Y(n845) );
  CLKBUFX2TS U1643 ( .A(n1511), .Y(n903) );
  CLKBUFX2TS U1644 ( .A(n903), .Y(n858) );
  CLKBUFX2TS U1645 ( .A(n843), .Y(n883) );
  CLKBUFX2TS U1646 ( .A(n883), .Y(n857) );
  AOI22X1TS U1647 ( .A0(n858), .A1(readOutBus[299]), .B0(n857), .B1(
        readOutBus[459]), .Y(n844) );
  NAND3XLTS U1648 ( .A(n846), .B(n845), .C(n844), .Y(readOut[139]) );
  AOI22X1TS U1649 ( .A0(n854), .A1(readOutBus[938]), .B0(n853), .B1(
        readOutBus[778]), .Y(n849) );
  AOI22X1TS U1650 ( .A0(n856), .A1(readOutBus[618]), .B0(n855), .B1(
        readOutBus[138]), .Y(n848) );
  AOI22X1TS U1651 ( .A0(n858), .A1(readOutBus[298]), .B0(n857), .B1(
        readOutBus[458]), .Y(n847) );
  NAND3XLTS U1652 ( .A(n849), .B(n848), .C(n847), .Y(readOut[138]) );
  AOI22X1TS U1653 ( .A0(n854), .A1(readOutBus[937]), .B0(n853), .B1(
        readOutBus[777]), .Y(n852) );
  AOI22X1TS U1654 ( .A0(n856), .A1(readOutBus[617]), .B0(n855), .B1(
        readOutBus[137]), .Y(n851) );
  AOI22X1TS U1655 ( .A0(n858), .A1(readOutBus[297]), .B0(n857), .B1(
        readOutBus[457]), .Y(n850) );
  NAND3XLTS U1656 ( .A(n852), .B(n851), .C(n850), .Y(readOut[137]) );
  AOI22X1TS U1657 ( .A0(n854), .A1(readOutBus[936]), .B0(n853), .B1(
        readOutBus[776]), .Y(n861) );
  AOI22X1TS U1658 ( .A0(n856), .A1(readOutBus[616]), .B0(n855), .B1(
        readOutBus[136]), .Y(n860) );
  AOI22X1TS U1659 ( .A0(n858), .A1(readOutBus[296]), .B0(n857), .B1(
        readOutBus[456]), .Y(n859) );
  NAND3XLTS U1660 ( .A(n861), .B(n860), .C(n859), .Y(readOut[136]) );
  CLKBUFX2TS U1661 ( .A(n880), .Y(n872) );
  CLKBUFX2TS U1662 ( .A(n881), .Y(n871) );
  AOI22X1TS U1663 ( .A0(n872), .A1(readOutBus[935]), .B0(n871), .B1(
        readOutBus[775]), .Y(n864) );
  CLKBUFX2TS U1664 ( .A(n902), .Y(n874) );
  CLKBUFX2TS U1665 ( .A(n882), .Y(n873) );
  AOI22X1TS U1666 ( .A0(n874), .A1(readOutBus[615]), .B0(n873), .B1(
        readOutBus[135]), .Y(n863) );
  CLKBUFX2TS U1667 ( .A(n903), .Y(n876) );
  CLKBUFX2TS U1668 ( .A(n883), .Y(n875) );
  AOI22X1TS U1669 ( .A0(n876), .A1(readOutBus[295]), .B0(n875), .B1(
        readOutBus[455]), .Y(n862) );
  NAND3XLTS U1670 ( .A(n864), .B(n863), .C(n862), .Y(readOut[135]) );
  AOI22X1TS U1671 ( .A0(n872), .A1(readOutBus[934]), .B0(n871), .B1(
        readOutBus[774]), .Y(n867) );
  AOI22X1TS U1672 ( .A0(n874), .A1(readOutBus[614]), .B0(n873), .B1(
        readOutBus[134]), .Y(n866) );
  AOI22X1TS U1673 ( .A0(n876), .A1(readOutBus[294]), .B0(n875), .B1(
        readOutBus[454]), .Y(n865) );
  NAND3XLTS U1674 ( .A(n867), .B(n866), .C(n865), .Y(readOut[134]) );
  AOI22X1TS U1675 ( .A0(n872), .A1(readOutBus[933]), .B0(n871), .B1(
        readOutBus[773]), .Y(n870) );
  AOI22X1TS U1676 ( .A0(n874), .A1(readOutBus[613]), .B0(n873), .B1(
        readOutBus[133]), .Y(n869) );
  AOI22X1TS U1677 ( .A0(n876), .A1(readOutBus[293]), .B0(n875), .B1(
        readOutBus[453]), .Y(n868) );
  NAND3XLTS U1678 ( .A(n870), .B(n869), .C(n868), .Y(readOut[133]) );
  AOI22X1TS U1679 ( .A0(n872), .A1(readOutBus[932]), .B0(n871), .B1(
        readOutBus[772]), .Y(n879) );
  AOI22X1TS U1680 ( .A0(n874), .A1(readOutBus[612]), .B0(n873), .B1(
        readOutBus[132]), .Y(n878) );
  AOI22X1TS U1681 ( .A0(n876), .A1(readOutBus[292]), .B0(n875), .B1(
        readOutBus[452]), .Y(n877) );
  NAND3XLTS U1682 ( .A(n879), .B(n878), .C(n877), .Y(readOut[132]) );
  CLKBUFX2TS U1683 ( .A(n880), .Y(n894) );
  CLKBUFX2TS U1684 ( .A(n881), .Y(n893) );
  AOI22X1TS U1685 ( .A0(n894), .A1(readOutBus[931]), .B0(n893), .B1(
        readOutBus[771]), .Y(n886) );
  CLKBUFX2TS U1686 ( .A(n902), .Y(n896) );
  CLKBUFX2TS U1687 ( .A(n882), .Y(n895) );
  AOI22X1TS U1688 ( .A0(n896), .A1(readOutBus[611]), .B0(n895), .B1(
        readOutBus[131]), .Y(n885) );
  CLKBUFX2TS U1689 ( .A(n903), .Y(n898) );
  CLKBUFX2TS U1690 ( .A(n883), .Y(n897) );
  AOI22X1TS U1691 ( .A0(n898), .A1(readOutBus[291]), .B0(n897), .B1(
        readOutBus[451]), .Y(n884) );
  NAND3XLTS U1692 ( .A(n886), .B(n885), .C(n884), .Y(readOut[131]) );
  AOI22X1TS U1693 ( .A0(n894), .A1(readOutBus[930]), .B0(n893), .B1(
        readOutBus[770]), .Y(n889) );
  AOI22X1TS U1694 ( .A0(n896), .A1(readOutBus[610]), .B0(n895), .B1(
        readOutBus[130]), .Y(n888) );
  AOI22X1TS U1695 ( .A0(n898), .A1(readOutBus[290]), .B0(n897), .B1(
        readOutBus[450]), .Y(n887) );
  NAND3XLTS U1696 ( .A(n889), .B(n888), .C(n887), .Y(readOut[130]) );
  AOI22X1TS U1697 ( .A0(n894), .A1(readOutBus[929]), .B0(n893), .B1(
        readOutBus[769]), .Y(n892) );
  AOI22X1TS U1698 ( .A0(n896), .A1(readOutBus[609]), .B0(n895), .B1(
        readOutBus[129]), .Y(n891) );
  AOI22X1TS U1699 ( .A0(n898), .A1(readOutBus[289]), .B0(n897), .B1(
        readOutBus[449]), .Y(n890) );
  NAND3XLTS U1700 ( .A(n892), .B(n891), .C(n890), .Y(readOut[129]) );
  AOI22X1TS U1701 ( .A0(n894), .A1(readOutBus[928]), .B0(n893), .B1(
        readOutBus[768]), .Y(n901) );
  AOI22X1TS U1702 ( .A0(n896), .A1(readOutBus[608]), .B0(n895), .B1(
        readOutBus[128]), .Y(n900) );
  AOI22X1TS U1703 ( .A0(n898), .A1(readOutBus[288]), .B0(n897), .B1(
        readOutBus[448]), .Y(n899) );
  NAND3XLTS U1704 ( .A(n901), .B(n900), .C(n899), .Y(readOut[128]) );
  CLKBUFX2TS U1705 ( .A(n1507), .Y(n1516) );
  CLKBUFX2TS U1706 ( .A(n1516), .Y(n914) );
  CLKBUFX2TS U1707 ( .A(n1506), .Y(n1417) );
  CLKBUFX2TS U1708 ( .A(n1417), .Y(n997) );
  CLKBUFX2TS U1709 ( .A(n997), .Y(n913) );
  AOI22X1TS U1710 ( .A0(n914), .A1(readOutBus[927]), .B0(n913), .B1(
        readOutBus[767]), .Y(n906) );
  CLKBUFX2TS U1711 ( .A(n902), .Y(n1418) );
  CLKBUFX2TS U1712 ( .A(n1418), .Y(n1478) );
  CLKBUFX2TS U1713 ( .A(n1478), .Y(n998) );
  CLKBUFX2TS U1714 ( .A(n998), .Y(n940) );
  CLKBUFX2TS U1715 ( .A(n940), .Y(n916) );
  CLKBUFX2TS U1716 ( .A(n1517), .Y(n999) );
  CLKBUFX2TS U1717 ( .A(n999), .Y(n915) );
  AOI22X1TS U1718 ( .A0(n916), .A1(readOutBus[607]), .B0(n915), .B1(
        readOutBus[127]), .Y(n905) );
  CLKBUFX2TS U1719 ( .A(n903), .Y(n1420) );
  CLKBUFX2TS U1720 ( .A(n1420), .Y(n1480) );
  CLKBUFX2TS U1721 ( .A(n1480), .Y(n1000) );
  CLKBUFX2TS U1722 ( .A(n1000), .Y(n941) );
  CLKBUFX2TS U1723 ( .A(n941), .Y(n918) );
  CLKBUFX2TS U1724 ( .A(n1519), .Y(n1001) );
  CLKBUFX2TS U1725 ( .A(n1001), .Y(n917) );
  AOI22X1TS U1726 ( .A0(n918), .A1(readOutBus[287]), .B0(n917), .B1(
        readOutBus[447]), .Y(n904) );
  NAND3XLTS U1727 ( .A(n906), .B(n905), .C(n904), .Y(readOut[127]) );
  AOI22X1TS U1728 ( .A0(n914), .A1(readOutBus[926]), .B0(n913), .B1(
        readOutBus[766]), .Y(n909) );
  AOI22X1TS U1729 ( .A0(n916), .A1(readOutBus[606]), .B0(n915), .B1(
        readOutBus[126]), .Y(n908) );
  AOI22X1TS U1730 ( .A0(n918), .A1(readOutBus[286]), .B0(n917), .B1(
        readOutBus[446]), .Y(n907) );
  NAND3XLTS U1731 ( .A(n909), .B(n908), .C(n907), .Y(readOut[126]) );
  AOI22X1TS U1732 ( .A0(n914), .A1(readOutBus[925]), .B0(n913), .B1(
        readOutBus[765]), .Y(n912) );
  AOI22X1TS U1733 ( .A0(n916), .A1(readOutBus[605]), .B0(n915), .B1(
        readOutBus[125]), .Y(n911) );
  AOI22X1TS U1734 ( .A0(n918), .A1(readOutBus[285]), .B0(n917), .B1(
        readOutBus[445]), .Y(n910) );
  NAND3XLTS U1735 ( .A(n912), .B(n911), .C(n910), .Y(readOut[125]) );
  AOI22X1TS U1736 ( .A0(n914), .A1(readOutBus[924]), .B0(n913), .B1(
        readOutBus[764]), .Y(n921) );
  AOI22X1TS U1737 ( .A0(n916), .A1(readOutBus[604]), .B0(n915), .B1(
        readOutBus[124]), .Y(n920) );
  AOI22X1TS U1738 ( .A0(n918), .A1(readOutBus[284]), .B0(n917), .B1(
        readOutBus[444]), .Y(n919) );
  NAND3XLTS U1739 ( .A(n921), .B(n920), .C(n919), .Y(readOut[124]) );
  CLKBUFX2TS U1740 ( .A(n1516), .Y(n932) );
  CLKBUFX2TS U1741 ( .A(n997), .Y(n931) );
  AOI22X1TS U1742 ( .A0(n932), .A1(readOutBus[923]), .B0(n931), .B1(
        readOutBus[763]), .Y(n924) );
  CLKBUFX2TS U1743 ( .A(n940), .Y(n934) );
  CLKBUFX2TS U1744 ( .A(n999), .Y(n933) );
  AOI22X1TS U1745 ( .A0(n934), .A1(readOutBus[603]), .B0(n933), .B1(
        readOutBus[123]), .Y(n923) );
  CLKBUFX2TS U1746 ( .A(n941), .Y(n936) );
  CLKBUFX2TS U1747 ( .A(n1001), .Y(n935) );
  AOI22X1TS U1748 ( .A0(n936), .A1(readOutBus[283]), .B0(n935), .B1(
        readOutBus[443]), .Y(n922) );
  NAND3XLTS U1749 ( .A(n924), .B(n923), .C(n922), .Y(readOut[123]) );
  AOI22X1TS U1750 ( .A0(n932), .A1(readOutBus[922]), .B0(n931), .B1(
        readOutBus[762]), .Y(n927) );
  AOI22X1TS U1751 ( .A0(n934), .A1(readOutBus[602]), .B0(n933), .B1(
        readOutBus[122]), .Y(n926) );
  AOI22X1TS U1752 ( .A0(n936), .A1(readOutBus[282]), .B0(n935), .B1(
        readOutBus[442]), .Y(n925) );
  NAND3XLTS U1753 ( .A(n927), .B(n926), .C(n925), .Y(readOut[122]) );
  AOI22X1TS U1754 ( .A0(n932), .A1(readOutBus[921]), .B0(n931), .B1(
        readOutBus[761]), .Y(n930) );
  AOI22X1TS U1755 ( .A0(n934), .A1(readOutBus[601]), .B0(n933), .B1(
        readOutBus[121]), .Y(n929) );
  AOI22X1TS U1756 ( .A0(n936), .A1(readOutBus[281]), .B0(n935), .B1(
        readOutBus[441]), .Y(n928) );
  NAND3XLTS U1757 ( .A(n930), .B(n929), .C(n928), .Y(readOut[121]) );
  AOI22X1TS U1758 ( .A0(n932), .A1(readOutBus[920]), .B0(n931), .B1(
        readOutBus[760]), .Y(n939) );
  AOI22X1TS U1759 ( .A0(n934), .A1(readOutBus[600]), .B0(n933), .B1(
        readOutBus[120]), .Y(n938) );
  AOI22X1TS U1760 ( .A0(n936), .A1(readOutBus[280]), .B0(n935), .B1(
        readOutBus[440]), .Y(n937) );
  NAND3XLTS U1761 ( .A(n939), .B(n938), .C(n937), .Y(readOut[120]) );
  CLKBUFX2TS U1762 ( .A(n1516), .Y(n952) );
  CLKBUFX2TS U1763 ( .A(n1080), .Y(n951) );
  AOI22X1TS U1764 ( .A0(n952), .A1(readOutBus[919]), .B0(n951), .B1(
        readOutBus[759]), .Y(n944) );
  CLKBUFX2TS U1765 ( .A(n940), .Y(n954) );
  CLKBUFX2TS U1766 ( .A(n1101), .Y(n953) );
  AOI22X1TS U1767 ( .A0(n954), .A1(readOutBus[599]), .B0(n953), .B1(
        readOutBus[119]), .Y(n943) );
  CLKBUFX2TS U1768 ( .A(n941), .Y(n956) );
  CLKBUFX2TS U1769 ( .A(n1102), .Y(n955) );
  AOI22X1TS U1770 ( .A0(n956), .A1(readOutBus[279]), .B0(n955), .B1(
        readOutBus[439]), .Y(n942) );
  NAND3XLTS U1771 ( .A(n944), .B(n943), .C(n942), .Y(readOut[119]) );
  AOI22X1TS U1772 ( .A0(n952), .A1(readOutBus[918]), .B0(n951), .B1(
        readOutBus[758]), .Y(n947) );
  AOI22X1TS U1773 ( .A0(n954), .A1(readOutBus[598]), .B0(n953), .B1(
        readOutBus[118]), .Y(n946) );
  AOI22X1TS U1774 ( .A0(n956), .A1(readOutBus[278]), .B0(n955), .B1(
        readOutBus[438]), .Y(n945) );
  NAND3XLTS U1775 ( .A(n947), .B(n946), .C(n945), .Y(readOut[118]) );
  AOI22X1TS U1776 ( .A0(n952), .A1(readOutBus[917]), .B0(n951), .B1(
        readOutBus[757]), .Y(n950) );
  AOI22X1TS U1777 ( .A0(n954), .A1(readOutBus[597]), .B0(n953), .B1(
        readOutBus[117]), .Y(n949) );
  AOI22X1TS U1778 ( .A0(n956), .A1(readOutBus[277]), .B0(n955), .B1(
        readOutBus[437]), .Y(n948) );
  NAND3XLTS U1779 ( .A(n950), .B(n949), .C(n948), .Y(readOut[117]) );
  AOI22X1TS U1780 ( .A0(n952), .A1(readOutBus[916]), .B0(n951), .B1(
        readOutBus[756]), .Y(n959) );
  AOI22X1TS U1781 ( .A0(n954), .A1(readOutBus[596]), .B0(n953), .B1(
        readOutBus[116]), .Y(n958) );
  AOI22X1TS U1782 ( .A0(n956), .A1(readOutBus[276]), .B0(n955), .B1(
        readOutBus[436]), .Y(n957) );
  NAND3XLTS U1783 ( .A(n959), .B(n958), .C(n957), .Y(readOut[116]) );
  CLKBUFX2TS U1784 ( .A(n1507), .Y(n1178) );
  CLKBUFX2TS U1785 ( .A(n1178), .Y(n1121) );
  CLKBUFX2TS U1786 ( .A(n1121), .Y(n1356) );
  CLKBUFX2TS U1787 ( .A(n1356), .Y(n1416) );
  CLKBUFX2TS U1788 ( .A(n1416), .Y(n1476) );
  CLKBUFX2TS U1789 ( .A(n1476), .Y(n996) );
  CLKBUFX2TS U1790 ( .A(n996), .Y(n970) );
  CLKBUFX2TS U1791 ( .A(n997), .Y(n969) );
  AOI22X1TS U1792 ( .A0(n970), .A1(readOutBus[915]), .B0(n969), .B1(
        readOutBus[755]), .Y(n962) );
  CLKBUFX2TS U1793 ( .A(n998), .Y(n972) );
  CLKBUFX2TS U1794 ( .A(n999), .Y(n971) );
  AOI22X1TS U1795 ( .A0(n972), .A1(readOutBus[595]), .B0(n971), .B1(
        readOutBus[115]), .Y(n961) );
  CLKBUFX2TS U1796 ( .A(n1000), .Y(n974) );
  CLKBUFX2TS U1797 ( .A(n1001), .Y(n973) );
  AOI22X1TS U1798 ( .A0(n974), .A1(readOutBus[275]), .B0(n973), .B1(
        readOutBus[435]), .Y(n960) );
  NAND3XLTS U1799 ( .A(n962), .B(n961), .C(n960), .Y(readOut[115]) );
  AOI22X1TS U1800 ( .A0(n970), .A1(readOutBus[914]), .B0(n969), .B1(
        readOutBus[754]), .Y(n965) );
  AOI22X1TS U1801 ( .A0(n972), .A1(readOutBus[594]), .B0(n971), .B1(
        readOutBus[114]), .Y(n964) );
  AOI22X1TS U1802 ( .A0(n974), .A1(readOutBus[274]), .B0(n973), .B1(
        readOutBus[434]), .Y(n963) );
  NAND3XLTS U1803 ( .A(n965), .B(n964), .C(n963), .Y(readOut[114]) );
  AOI22X1TS U1804 ( .A0(n970), .A1(readOutBus[913]), .B0(n969), .B1(
        readOutBus[753]), .Y(n968) );
  AOI22X1TS U1805 ( .A0(n972), .A1(readOutBus[593]), .B0(n971), .B1(
        readOutBus[113]), .Y(n967) );
  AOI22X1TS U1806 ( .A0(n974), .A1(readOutBus[273]), .B0(n973), .B1(
        readOutBus[433]), .Y(n966) );
  NAND3XLTS U1807 ( .A(n968), .B(n967), .C(n966), .Y(readOut[113]) );
  AOI22X1TS U1808 ( .A0(n970), .A1(readOutBus[912]), .B0(n969), .B1(
        readOutBus[752]), .Y(n977) );
  AOI22X1TS U1809 ( .A0(n972), .A1(readOutBus[592]), .B0(n971), .B1(
        readOutBus[112]), .Y(n976) );
  AOI22X1TS U1810 ( .A0(n974), .A1(readOutBus[272]), .B0(n973), .B1(
        readOutBus[432]), .Y(n975) );
  NAND3XLTS U1811 ( .A(n977), .B(n976), .C(n975), .Y(readOut[112]) );
  CLKBUFX2TS U1812 ( .A(n996), .Y(n988) );
  CLKBUFX2TS U1813 ( .A(n1080), .Y(n1357) );
  CLKBUFX2TS U1814 ( .A(n1357), .Y(n987) );
  AOI22X1TS U1815 ( .A0(n988), .A1(readOutBus[911]), .B0(n987), .B1(
        readOutBus[751]), .Y(n980) );
  CLKBUFX2TS U1816 ( .A(n998), .Y(n1058) );
  CLKBUFX2TS U1817 ( .A(n1058), .Y(n990) );
  CLKBUFX2TS U1818 ( .A(n1101), .Y(n1359) );
  CLKBUFX2TS U1819 ( .A(n1359), .Y(n989) );
  AOI22X1TS U1820 ( .A0(n990), .A1(readOutBus[591]), .B0(n989), .B1(
        readOutBus[111]), .Y(n979) );
  CLKBUFX2TS U1821 ( .A(n1000), .Y(n1060) );
  CLKBUFX2TS U1822 ( .A(n1060), .Y(n992) );
  CLKBUFX2TS U1823 ( .A(n1102), .Y(n1361) );
  CLKBUFX2TS U1824 ( .A(n1361), .Y(n991) );
  AOI22X1TS U1825 ( .A0(n992), .A1(readOutBus[271]), .B0(n991), .B1(
        readOutBus[431]), .Y(n978) );
  NAND3XLTS U1826 ( .A(n980), .B(n979), .C(n978), .Y(readOut[111]) );
  AOI22X1TS U1827 ( .A0(n988), .A1(readOutBus[910]), .B0(n987), .B1(
        readOutBus[750]), .Y(n983) );
  AOI22X1TS U1828 ( .A0(n990), .A1(readOutBus[590]), .B0(n989), .B1(
        readOutBus[110]), .Y(n982) );
  AOI22X1TS U1829 ( .A0(n992), .A1(readOutBus[270]), .B0(n991), .B1(
        readOutBus[430]), .Y(n981) );
  NAND3XLTS U1830 ( .A(n983), .B(n982), .C(n981), .Y(readOut[110]) );
  AOI22X1TS U1831 ( .A0(n988), .A1(readOutBus[909]), .B0(n987), .B1(
        readOutBus[749]), .Y(n986) );
  AOI22X1TS U1832 ( .A0(n990), .A1(readOutBus[589]), .B0(n989), .B1(
        readOutBus[109]), .Y(n985) );
  AOI22X1TS U1833 ( .A0(n992), .A1(readOutBus[269]), .B0(n991), .B1(
        readOutBus[429]), .Y(n984) );
  NAND3XLTS U1834 ( .A(n986), .B(n985), .C(n984), .Y(readOut[109]) );
  AOI22X1TS U1835 ( .A0(n988), .A1(readOutBus[908]), .B0(n987), .B1(
        readOutBus[748]), .Y(n995) );
  AOI22X1TS U1836 ( .A0(n990), .A1(readOutBus[588]), .B0(n989), .B1(
        readOutBus[108]), .Y(n994) );
  AOI22X1TS U1837 ( .A0(n992), .A1(readOutBus[268]), .B0(n991), .B1(
        readOutBus[428]), .Y(n993) );
  NAND3XLTS U1838 ( .A(n995), .B(n994), .C(n993), .Y(readOut[108]) );
  CLKBUFX2TS U1839 ( .A(n996), .Y(n1012) );
  CLKBUFX2TS U1840 ( .A(n997), .Y(n1057) );
  CLKBUFX2TS U1841 ( .A(n1057), .Y(n1011) );
  AOI22X1TS U1842 ( .A0(n1012), .A1(readOutBus[907]), .B0(n1011), .B1(
        readOutBus[747]), .Y(n1004) );
  CLKBUFX2TS U1843 ( .A(n998), .Y(n1014) );
  CLKBUFX2TS U1844 ( .A(n999), .Y(n1059) );
  CLKBUFX2TS U1845 ( .A(n1059), .Y(n1013) );
  AOI22X1TS U1846 ( .A0(n1014), .A1(readOutBus[587]), .B0(n1013), .B1(
        readOutBus[107]), .Y(n1003) );
  CLKBUFX2TS U1847 ( .A(n1000), .Y(n1016) );
  CLKBUFX2TS U1848 ( .A(n1001), .Y(n1061) );
  CLKBUFX2TS U1849 ( .A(n1061), .Y(n1015) );
  AOI22X1TS U1850 ( .A0(n1016), .A1(readOutBus[267]), .B0(n1015), .B1(
        readOutBus[427]), .Y(n1002) );
  NAND3XLTS U1851 ( .A(n1004), .B(n1003), .C(n1002), .Y(readOut[107]) );
  AOI22X1TS U1852 ( .A0(n1012), .A1(readOutBus[906]), .B0(n1011), .B1(
        readOutBus[746]), .Y(n1007) );
  AOI22X1TS U1853 ( .A0(n1014), .A1(readOutBus[586]), .B0(n1013), .B1(
        readOutBus[106]), .Y(n1006) );
  AOI22X1TS U1854 ( .A0(n1016), .A1(readOutBus[266]), .B0(n1015), .B1(
        readOutBus[426]), .Y(n1005) );
  NAND3XLTS U1855 ( .A(n1007), .B(n1006), .C(n1005), .Y(readOut[106]) );
  AOI22X1TS U1856 ( .A0(n1012), .A1(readOutBus[905]), .B0(n1011), .B1(
        readOutBus[745]), .Y(n1010) );
  AOI22X1TS U1857 ( .A0(n1014), .A1(readOutBus[585]), .B0(n1013), .B1(
        readOutBus[105]), .Y(n1009) );
  AOI22X1TS U1858 ( .A0(n1016), .A1(readOutBus[265]), .B0(n1015), .B1(
        readOutBus[425]), .Y(n1008) );
  NAND3XLTS U1859 ( .A(n1010), .B(n1009), .C(n1008), .Y(readOut[105]) );
  AOI22X1TS U1860 ( .A0(n1012), .A1(readOutBus[904]), .B0(n1011), .B1(
        readOutBus[744]), .Y(n1019) );
  AOI22X1TS U1861 ( .A0(n1014), .A1(readOutBus[584]), .B0(n1013), .B1(
        readOutBus[104]), .Y(n1018) );
  AOI22X1TS U1862 ( .A0(n1016), .A1(readOutBus[264]), .B0(n1015), .B1(
        readOutBus[424]), .Y(n1017) );
  NAND3XLTS U1863 ( .A(n1019), .B(n1018), .C(n1017), .Y(readOut[104]) );
  CLKBUFX2TS U1864 ( .A(n1056), .Y(n1030) );
  CLKBUFX2TS U1865 ( .A(n1057), .Y(n1029) );
  AOI22X1TS U1866 ( .A0(n1030), .A1(readOutBus[903]), .B0(n1029), .B1(
        readOutBus[743]), .Y(n1022) );
  CLKBUFX2TS U1867 ( .A(n1058), .Y(n1032) );
  CLKBUFX2TS U1868 ( .A(n1059), .Y(n1031) );
  AOI22X1TS U1869 ( .A0(n1032), .A1(readOutBus[583]), .B0(n1031), .B1(
        readOutBus[103]), .Y(n1021) );
  CLKBUFX2TS U1870 ( .A(n1060), .Y(n1034) );
  CLKBUFX2TS U1871 ( .A(n1061), .Y(n1033) );
  AOI22X1TS U1872 ( .A0(n1034), .A1(readOutBus[263]), .B0(n1033), .B1(
        readOutBus[423]), .Y(n1020) );
  NAND3XLTS U1873 ( .A(n1022), .B(n1021), .C(n1020), .Y(readOut[103]) );
  AOI22X1TS U1874 ( .A0(n1030), .A1(readOutBus[902]), .B0(n1029), .B1(
        readOutBus[742]), .Y(n1025) );
  AOI22X1TS U1875 ( .A0(n1032), .A1(readOutBus[582]), .B0(n1031), .B1(
        readOutBus[102]), .Y(n1024) );
  AOI22X1TS U1876 ( .A0(n1034), .A1(readOutBus[262]), .B0(n1033), .B1(
        readOutBus[422]), .Y(n1023) );
  NAND3XLTS U1877 ( .A(n1025), .B(n1024), .C(n1023), .Y(readOut[102]) );
  AOI22X1TS U1878 ( .A0(n1030), .A1(readOutBus[901]), .B0(n1029), .B1(
        readOutBus[741]), .Y(n1028) );
  AOI22X1TS U1879 ( .A0(n1032), .A1(readOutBus[581]), .B0(n1031), .B1(
        readOutBus[101]), .Y(n1027) );
  AOI22X1TS U1880 ( .A0(n1034), .A1(readOutBus[261]), .B0(n1033), .B1(
        readOutBus[421]), .Y(n1026) );
  NAND3XLTS U1881 ( .A(n1028), .B(n1027), .C(n1026), .Y(readOut[101]) );
  AOI22X1TS U1882 ( .A0(n1030), .A1(readOutBus[900]), .B0(n1029), .B1(
        readOutBus[740]), .Y(n1037) );
  AOI22X1TS U1883 ( .A0(n1032), .A1(readOutBus[580]), .B0(n1031), .B1(
        readOutBus[100]), .Y(n1036) );
  AOI22X1TS U1884 ( .A0(n1034), .A1(readOutBus[260]), .B0(n1033), .B1(
        readOutBus[420]), .Y(n1035) );
  NAND3XLTS U1885 ( .A(n1037), .B(n1036), .C(n1035), .Y(readOut[100]) );
  CLKBUFX2TS U1886 ( .A(n1056), .Y(n1048) );
  CLKBUFX2TS U1887 ( .A(n1057), .Y(n1047) );
  AOI22X1TS U1888 ( .A0(n1048), .A1(readOutBus[899]), .B0(n1047), .B1(
        readOutBus[739]), .Y(n1040) );
  CLKBUFX2TS U1889 ( .A(n1058), .Y(n1050) );
  CLKBUFX2TS U1890 ( .A(n1059), .Y(n1049) );
  AOI22X1TS U1891 ( .A0(n1050), .A1(readOutBus[579]), .B0(n1049), .B1(
        readOutBus[99]), .Y(n1039) );
  CLKBUFX2TS U1892 ( .A(n1060), .Y(n1052) );
  CLKBUFX2TS U1893 ( .A(n1061), .Y(n1051) );
  AOI22X1TS U1894 ( .A0(n1052), .A1(readOutBus[259]), .B0(n1051), .B1(
        readOutBus[419]), .Y(n1038) );
  NAND3XLTS U1895 ( .A(n1040), .B(n1039), .C(n1038), .Y(readOut[99]) );
  AOI22X1TS U1896 ( .A0(n1048), .A1(readOutBus[898]), .B0(n1047), .B1(
        readOutBus[738]), .Y(n1043) );
  AOI22X1TS U1897 ( .A0(n1050), .A1(readOutBus[578]), .B0(n1049), .B1(
        readOutBus[98]), .Y(n1042) );
  AOI22X1TS U1898 ( .A0(n1052), .A1(readOutBus[258]), .B0(n1051), .B1(
        readOutBus[418]), .Y(n1041) );
  NAND3XLTS U1899 ( .A(n1043), .B(n1042), .C(n1041), .Y(readOut[98]) );
  AOI22X1TS U1900 ( .A0(n1048), .A1(readOutBus[897]), .B0(n1047), .B1(
        readOutBus[737]), .Y(n1046) );
  AOI22X1TS U1901 ( .A0(n1050), .A1(readOutBus[577]), .B0(n1049), .B1(
        readOutBus[97]), .Y(n1045) );
  AOI22X1TS U1902 ( .A0(n1052), .A1(readOutBus[257]), .B0(n1051), .B1(
        readOutBus[417]), .Y(n1044) );
  NAND3XLTS U1903 ( .A(n1046), .B(n1045), .C(n1044), .Y(readOut[97]) );
  AOI22X1TS U1904 ( .A0(n1048), .A1(readOutBus[896]), .B0(n1047), .B1(
        readOutBus[736]), .Y(n1055) );
  AOI22X1TS U1905 ( .A0(n1050), .A1(readOutBus[576]), .B0(n1049), .B1(
        readOutBus[96]), .Y(n1054) );
  AOI22X1TS U1906 ( .A0(n1052), .A1(readOutBus[256]), .B0(n1051), .B1(
        readOutBus[416]), .Y(n1053) );
  NAND3XLTS U1907 ( .A(n1055), .B(n1054), .C(n1053), .Y(readOut[96]) );
  CLKBUFX2TS U1908 ( .A(n1056), .Y(n1072) );
  CLKBUFX2TS U1909 ( .A(n1057), .Y(n1071) );
  AOI22X1TS U1910 ( .A0(n1072), .A1(readOutBus[895]), .B0(n1071), .B1(
        readOutBus[735]), .Y(n1064) );
  CLKBUFX2TS U1911 ( .A(n1058), .Y(n1074) );
  CLKBUFX2TS U1912 ( .A(n1059), .Y(n1073) );
  AOI22X1TS U1913 ( .A0(n1074), .A1(readOutBus[575]), .B0(n1073), .B1(
        readOutBus[95]), .Y(n1063) );
  CLKBUFX2TS U1914 ( .A(n1060), .Y(n1076) );
  CLKBUFX2TS U1915 ( .A(n1061), .Y(n1075) );
  AOI22X1TS U1916 ( .A0(n1076), .A1(readOutBus[255]), .B0(n1075), .B1(
        readOutBus[415]), .Y(n1062) );
  NAND3XLTS U1917 ( .A(n1064), .B(n1063), .C(n1062), .Y(readOut[95]) );
  AOI22X1TS U1918 ( .A0(n1072), .A1(readOutBus[894]), .B0(n1071), .B1(
        readOutBus[734]), .Y(n1067) );
  AOI22X1TS U1919 ( .A0(n1074), .A1(readOutBus[574]), .B0(n1073), .B1(
        readOutBus[94]), .Y(n1066) );
  AOI22X1TS U1920 ( .A0(n1076), .A1(readOutBus[254]), .B0(n1075), .B1(
        readOutBus[414]), .Y(n1065) );
  NAND3XLTS U1921 ( .A(n1067), .B(n1066), .C(n1065), .Y(readOut[94]) );
  AOI22X1TS U1922 ( .A0(n1072), .A1(readOutBus[893]), .B0(n1071), .B1(
        readOutBus[733]), .Y(n1070) );
  AOI22X1TS U1923 ( .A0(n1074), .A1(readOutBus[573]), .B0(n1073), .B1(
        readOutBus[93]), .Y(n1069) );
  AOI22X1TS U1924 ( .A0(n1076), .A1(readOutBus[253]), .B0(n1075), .B1(
        readOutBus[413]), .Y(n1068) );
  NAND3XLTS U1925 ( .A(n1070), .B(n1069), .C(n1068), .Y(readOut[93]) );
  AOI22X1TS U1926 ( .A0(n1072), .A1(readOutBus[892]), .B0(n1071), .B1(
        readOutBus[732]), .Y(n1079) );
  AOI22X1TS U1927 ( .A0(n1074), .A1(readOutBus[572]), .B0(n1073), .B1(
        readOutBus[92]), .Y(n1078) );
  AOI22X1TS U1928 ( .A0(n1076), .A1(readOutBus[252]), .B0(n1075), .B1(
        readOutBus[412]), .Y(n1077) );
  NAND3XLTS U1929 ( .A(n1079), .B(n1078), .C(n1077), .Y(readOut[92]) );
  CLKBUFX2TS U1930 ( .A(n1121), .Y(n1093) );
  CLKBUFX2TS U1931 ( .A(n1080), .Y(n1515) );
  CLKBUFX2TS U1932 ( .A(n1515), .Y(n1092) );
  AOI22X1TS U1933 ( .A0(n1093), .A1(readOutBus[891]), .B0(n1092), .B1(
        readOutBus[731]), .Y(n1085) );
  CLKBUFX2TS U1934 ( .A(n1081), .Y(n1180) );
  CLKBUFX2TS U1935 ( .A(n1180), .Y(n1122) );
  CLKBUFX2TS U1936 ( .A(n1122), .Y(n1095) );
  CLKBUFX2TS U1937 ( .A(n1517), .Y(n1094) );
  AOI22X1TS U1938 ( .A0(n1095), .A1(readOutBus[571]), .B0(n1094), .B1(
        readOutBus[91]), .Y(n1084) );
  CLKBUFX2TS U1939 ( .A(n1082), .Y(n1182) );
  CLKBUFX2TS U1940 ( .A(n1182), .Y(n1123) );
  CLKBUFX2TS U1941 ( .A(n1123), .Y(n1097) );
  CLKBUFX2TS U1942 ( .A(n1519), .Y(n1096) );
  AOI22X1TS U1943 ( .A0(n1097), .A1(readOutBus[251]), .B0(n1096), .B1(
        readOutBus[411]), .Y(n1083) );
  NAND3XLTS U1944 ( .A(n1085), .B(n1084), .C(n1083), .Y(readOut[91]) );
  AOI22X1TS U1945 ( .A0(n1093), .A1(readOutBus[890]), .B0(n1092), .B1(
        readOutBus[730]), .Y(n1088) );
  AOI22X1TS U1946 ( .A0(n1095), .A1(readOutBus[570]), .B0(n1094), .B1(
        readOutBus[90]), .Y(n1087) );
  AOI22X1TS U1947 ( .A0(n1097), .A1(readOutBus[250]), .B0(n1096), .B1(
        readOutBus[410]), .Y(n1086) );
  NAND3XLTS U1948 ( .A(n1088), .B(n1087), .C(n1086), .Y(readOut[90]) );
  AOI22X1TS U1949 ( .A0(n1093), .A1(readOutBus[889]), .B0(n1092), .B1(
        readOutBus[729]), .Y(n1091) );
  AOI22X1TS U1950 ( .A0(n1095), .A1(readOutBus[569]), .B0(n1094), .B1(
        readOutBus[89]), .Y(n1090) );
  AOI22X1TS U1951 ( .A0(n1097), .A1(readOutBus[249]), .B0(n1096), .B1(
        readOutBus[409]), .Y(n1089) );
  NAND3XLTS U1952 ( .A(n1091), .B(n1090), .C(n1089), .Y(readOut[89]) );
  AOI22X1TS U1953 ( .A0(n1093), .A1(readOutBus[888]), .B0(n1092), .B1(
        readOutBus[728]), .Y(n1100) );
  AOI22X1TS U1954 ( .A0(n1095), .A1(readOutBus[568]), .B0(n1094), .B1(
        readOutBus[88]), .Y(n1099) );
  AOI22X1TS U1955 ( .A0(n1097), .A1(readOutBus[248]), .B0(n1096), .B1(
        readOutBus[408]), .Y(n1098) );
  NAND3XLTS U1956 ( .A(n1100), .B(n1099), .C(n1098), .Y(readOut[88]) );
  CLKBUFX2TS U1957 ( .A(n1121), .Y(n1113) );
  CLKBUFX2TS U1958 ( .A(n1515), .Y(n1112) );
  AOI22X1TS U1959 ( .A0(n1113), .A1(readOutBus[887]), .B0(n1112), .B1(
        readOutBus[727]), .Y(n1105) );
  CLKBUFX2TS U1960 ( .A(n1122), .Y(n1115) );
  CLKBUFX2TS U1961 ( .A(n1101), .Y(n1114) );
  AOI22X1TS U1962 ( .A0(n1115), .A1(readOutBus[567]), .B0(n1114), .B1(
        readOutBus[87]), .Y(n1104) );
  CLKBUFX2TS U1963 ( .A(n1123), .Y(n1117) );
  CLKBUFX2TS U1964 ( .A(n1102), .Y(n1116) );
  AOI22X1TS U1965 ( .A0(n1117), .A1(readOutBus[247]), .B0(n1116), .B1(
        readOutBus[407]), .Y(n1103) );
  NAND3XLTS U1966 ( .A(n1105), .B(n1104), .C(n1103), .Y(readOut[87]) );
  AOI22X1TS U1967 ( .A0(n1113), .A1(readOutBus[886]), .B0(n1112), .B1(
        readOutBus[726]), .Y(n1108) );
  AOI22X1TS U1968 ( .A0(n1115), .A1(readOutBus[566]), .B0(n1114), .B1(
        readOutBus[86]), .Y(n1107) );
  AOI22X1TS U1969 ( .A0(n1117), .A1(readOutBus[246]), .B0(n1116), .B1(
        readOutBus[406]), .Y(n1106) );
  NAND3XLTS U1970 ( .A(n1108), .B(n1107), .C(n1106), .Y(readOut[86]) );
  AOI22X1TS U1971 ( .A0(n1113), .A1(readOutBus[885]), .B0(n1112), .B1(
        readOutBus[725]), .Y(n1111) );
  AOI22X1TS U1972 ( .A0(n1115), .A1(readOutBus[565]), .B0(n1114), .B1(
        readOutBus[85]), .Y(n1110) );
  AOI22X1TS U1973 ( .A0(n1117), .A1(readOutBus[245]), .B0(n1116), .B1(
        readOutBus[405]), .Y(n1109) );
  NAND3XLTS U1974 ( .A(n1111), .B(n1110), .C(n1109), .Y(readOut[85]) );
  AOI22X1TS U1975 ( .A0(n1113), .A1(readOutBus[884]), .B0(n1112), .B1(
        readOutBus[724]), .Y(n1120) );
  AOI22X1TS U1976 ( .A0(n1115), .A1(readOutBus[564]), .B0(n1114), .B1(
        readOutBus[84]), .Y(n1119) );
  AOI22X1TS U1977 ( .A0(n1117), .A1(readOutBus[244]), .B0(n1116), .B1(
        readOutBus[404]), .Y(n1118) );
  NAND3XLTS U1978 ( .A(n1120), .B(n1119), .C(n1118), .Y(readOut[84]) );
  CLKBUFX2TS U1979 ( .A(n1121), .Y(n1134) );
  CLKBUFX2TS U1980 ( .A(n1515), .Y(n1133) );
  AOI22X1TS U1981 ( .A0(n1134), .A1(readOutBus[883]), .B0(n1133), .B1(
        readOutBus[723]), .Y(n1126) );
  CLKBUFX2TS U1982 ( .A(n1122), .Y(n1136) );
  CLKBUFX2TS U1983 ( .A(n1508), .Y(n1419) );
  CLKBUFX2TS U1984 ( .A(n1419), .Y(n1135) );
  AOI22X1TS U1985 ( .A0(n1136), .A1(readOutBus[563]), .B0(n1135), .B1(
        readOutBus[83]), .Y(n1125) );
  CLKBUFX2TS U1986 ( .A(n1123), .Y(n1138) );
  CLKBUFX2TS U1987 ( .A(n1510), .Y(n1421) );
  CLKBUFX2TS U1988 ( .A(n1421), .Y(n1137) );
  AOI22X1TS U1989 ( .A0(n1138), .A1(readOutBus[243]), .B0(n1137), .B1(
        readOutBus[403]), .Y(n1124) );
  NAND3XLTS U1990 ( .A(n1126), .B(n1125), .C(n1124), .Y(readOut[83]) );
  AOI22X1TS U1991 ( .A0(n1134), .A1(readOutBus[882]), .B0(n1133), .B1(
        readOutBus[722]), .Y(n1129) );
  AOI22X1TS U1992 ( .A0(n1136), .A1(readOutBus[562]), .B0(n1135), .B1(
        readOutBus[82]), .Y(n1128) );
  AOI22X1TS U1993 ( .A0(n1138), .A1(readOutBus[242]), .B0(n1137), .B1(
        readOutBus[402]), .Y(n1127) );
  NAND3XLTS U1994 ( .A(n1129), .B(n1128), .C(n1127), .Y(readOut[82]) );
  AOI22X1TS U1995 ( .A0(n1134), .A1(readOutBus[881]), .B0(n1133), .B1(
        readOutBus[721]), .Y(n1132) );
  AOI22X1TS U1996 ( .A0(n1136), .A1(readOutBus[561]), .B0(n1135), .B1(
        readOutBus[81]), .Y(n1131) );
  AOI22X1TS U1997 ( .A0(n1138), .A1(readOutBus[241]), .B0(n1137), .B1(
        readOutBus[401]), .Y(n1130) );
  NAND3XLTS U1998 ( .A(n1132), .B(n1131), .C(n1130), .Y(readOut[81]) );
  AOI22X1TS U1999 ( .A0(n1134), .A1(readOutBus[880]), .B0(n1133), .B1(
        readOutBus[720]), .Y(n1141) );
  AOI22X1TS U2000 ( .A0(n1136), .A1(readOutBus[560]), .B0(n1135), .B1(
        readOutBus[80]), .Y(n1140) );
  AOI22X1TS U2001 ( .A0(n1138), .A1(readOutBus[240]), .B0(n1137), .B1(
        readOutBus[400]), .Y(n1139) );
  NAND3XLTS U2002 ( .A(n1141), .B(n1140), .C(n1139), .Y(readOut[80]) );
  CLKBUFX2TS U2003 ( .A(n1178), .Y(n1152) );
  CLKBUFX2TS U2004 ( .A(n1179), .Y(n1151) );
  AOI22X1TS U2005 ( .A0(n1152), .A1(readOutBus[879]), .B0(n1151), .B1(
        readOutBus[719]), .Y(n1144) );
  CLKBUFX2TS U2006 ( .A(n1180), .Y(n1154) );
  CLKBUFX2TS U2007 ( .A(n1181), .Y(n1153) );
  AOI22X1TS U2008 ( .A0(n1154), .A1(readOutBus[559]), .B0(n1153), .B1(
        readOutBus[79]), .Y(n1143) );
  CLKBUFX2TS U2009 ( .A(n1182), .Y(n1156) );
  CLKBUFX2TS U2010 ( .A(n1183), .Y(n1155) );
  AOI22X1TS U2011 ( .A0(n1156), .A1(readOutBus[239]), .B0(n1155), .B1(
        readOutBus[399]), .Y(n1142) );
  NAND3XLTS U2012 ( .A(n1144), .B(n1143), .C(n1142), .Y(readOut[79]) );
  AOI22X1TS U2013 ( .A0(n1152), .A1(readOutBus[878]), .B0(n1151), .B1(
        readOutBus[718]), .Y(n1147) );
  AOI22X1TS U2014 ( .A0(n1154), .A1(readOutBus[558]), .B0(n1153), .B1(
        readOutBus[78]), .Y(n1146) );
  AOI22X1TS U2015 ( .A0(n1156), .A1(readOutBus[238]), .B0(n1155), .B1(
        readOutBus[398]), .Y(n1145) );
  NAND3XLTS U2016 ( .A(n1147), .B(n1146), .C(n1145), .Y(readOut[78]) );
  AOI22X1TS U2017 ( .A0(n1152), .A1(readOutBus[877]), .B0(n1151), .B1(
        readOutBus[717]), .Y(n1150) );
  AOI22X1TS U2018 ( .A0(n1154), .A1(readOutBus[557]), .B0(n1153), .B1(
        readOutBus[77]), .Y(n1149) );
  AOI22X1TS U2019 ( .A0(n1156), .A1(readOutBus[237]), .B0(n1155), .B1(
        readOutBus[397]), .Y(n1148) );
  NAND3XLTS U2020 ( .A(n1150), .B(n1149), .C(n1148), .Y(readOut[77]) );
  AOI22X1TS U2021 ( .A0(n1152), .A1(readOutBus[876]), .B0(n1151), .B1(
        readOutBus[716]), .Y(n1159) );
  AOI22X1TS U2022 ( .A0(n1154), .A1(readOutBus[556]), .B0(n1153), .B1(
        readOutBus[76]), .Y(n1158) );
  AOI22X1TS U2023 ( .A0(n1156), .A1(readOutBus[236]), .B0(n1155), .B1(
        readOutBus[396]), .Y(n1157) );
  NAND3XLTS U2024 ( .A(n1159), .B(n1158), .C(n1157), .Y(readOut[76]) );
  CLKBUFX2TS U2025 ( .A(n1178), .Y(n1238) );
  CLKBUFX2TS U2026 ( .A(n1238), .Y(n1170) );
  CLKBUFX2TS U2027 ( .A(n1179), .Y(n1169) );
  AOI22X1TS U2028 ( .A0(n1170), .A1(readOutBus[875]), .B0(n1169), .B1(
        readOutBus[715]), .Y(n1162) );
  CLKBUFX2TS U2029 ( .A(n1180), .Y(n1240) );
  CLKBUFX2TS U2030 ( .A(n1240), .Y(n1172) );
  CLKBUFX2TS U2031 ( .A(n1181), .Y(n1171) );
  AOI22X1TS U2032 ( .A0(n1172), .A1(readOutBus[555]), .B0(n1171), .B1(
        readOutBus[75]), .Y(n1161) );
  CLKBUFX2TS U2033 ( .A(n1182), .Y(n1242) );
  CLKBUFX2TS U2034 ( .A(n1242), .Y(n1174) );
  CLKBUFX2TS U2035 ( .A(n1183), .Y(n1173) );
  AOI22X1TS U2036 ( .A0(n1174), .A1(readOutBus[235]), .B0(n1173), .B1(
        readOutBus[395]), .Y(n1160) );
  NAND3XLTS U2037 ( .A(n1162), .B(n1161), .C(n1160), .Y(readOut[75]) );
  AOI22X1TS U2038 ( .A0(n1170), .A1(readOutBus[874]), .B0(n1169), .B1(
        readOutBus[714]), .Y(n1165) );
  AOI22X1TS U2039 ( .A0(n1172), .A1(readOutBus[554]), .B0(n1171), .B1(
        readOutBus[74]), .Y(n1164) );
  AOI22X1TS U2040 ( .A0(n1174), .A1(readOutBus[234]), .B0(n1173), .B1(
        readOutBus[394]), .Y(n1163) );
  NAND3XLTS U2041 ( .A(n1165), .B(n1164), .C(n1163), .Y(readOut[74]) );
  AOI22X1TS U2042 ( .A0(n1170), .A1(readOutBus[873]), .B0(n1169), .B1(
        readOutBus[713]), .Y(n1168) );
  AOI22X1TS U2043 ( .A0(n1172), .A1(readOutBus[553]), .B0(n1171), .B1(
        readOutBus[73]), .Y(n1167) );
  AOI22X1TS U2044 ( .A0(n1174), .A1(readOutBus[233]), .B0(n1173), .B1(
        readOutBus[393]), .Y(n1166) );
  NAND3XLTS U2045 ( .A(n1168), .B(n1167), .C(n1166), .Y(readOut[73]) );
  AOI22X1TS U2046 ( .A0(n1170), .A1(readOutBus[872]), .B0(n1169), .B1(
        readOutBus[712]), .Y(n1177) );
  AOI22X1TS U2047 ( .A0(n1172), .A1(readOutBus[552]), .B0(n1171), .B1(
        readOutBus[72]), .Y(n1176) );
  AOI22X1TS U2048 ( .A0(n1174), .A1(readOutBus[232]), .B0(n1173), .B1(
        readOutBus[392]), .Y(n1175) );
  NAND3XLTS U2049 ( .A(n1177), .B(n1176), .C(n1175), .Y(readOut[72]) );
  CLKBUFX2TS U2050 ( .A(n1178), .Y(n1194) );
  CLKBUFX2TS U2051 ( .A(n1179), .Y(n1193) );
  AOI22X1TS U2052 ( .A0(n1194), .A1(readOutBus[871]), .B0(n1193), .B1(
        readOutBus[711]), .Y(n1186) );
  CLKBUFX2TS U2053 ( .A(n1180), .Y(n1196) );
  CLKBUFX2TS U2054 ( .A(n1181), .Y(n1195) );
  AOI22X1TS U2055 ( .A0(n1196), .A1(readOutBus[551]), .B0(n1195), .B1(
        readOutBus[71]), .Y(n1185) );
  CLKBUFX2TS U2056 ( .A(n1182), .Y(n1198) );
  CLKBUFX2TS U2057 ( .A(n1183), .Y(n1197) );
  AOI22X1TS U2058 ( .A0(n1198), .A1(readOutBus[231]), .B0(n1197), .B1(
        readOutBus[391]), .Y(n1184) );
  NAND3XLTS U2059 ( .A(n1186), .B(n1185), .C(n1184), .Y(readOut[71]) );
  AOI22X1TS U2060 ( .A0(n1194), .A1(readOutBus[870]), .B0(n1193), .B1(
        readOutBus[710]), .Y(n1189) );
  AOI22X1TS U2061 ( .A0(n1196), .A1(readOutBus[550]), .B0(n1195), .B1(
        readOutBus[70]), .Y(n1188) );
  AOI22X1TS U2062 ( .A0(n1198), .A1(readOutBus[230]), .B0(n1197), .B1(
        readOutBus[390]), .Y(n1187) );
  NAND3XLTS U2063 ( .A(n1189), .B(n1188), .C(n1187), .Y(readOut[70]) );
  AOI22X1TS U2064 ( .A0(n1194), .A1(readOutBus[869]), .B0(n1193), .B1(
        readOutBus[709]), .Y(n1192) );
  AOI22X1TS U2065 ( .A0(n1196), .A1(readOutBus[549]), .B0(n1195), .B1(
        readOutBus[69]), .Y(n1191) );
  AOI22X1TS U2066 ( .A0(n1198), .A1(readOutBus[229]), .B0(n1197), .B1(
        readOutBus[389]), .Y(n1190) );
  NAND3XLTS U2067 ( .A(n1192), .B(n1191), .C(n1190), .Y(readOut[69]) );
  AOI22X1TS U2068 ( .A0(n1194), .A1(readOutBus[868]), .B0(n1193), .B1(
        readOutBus[708]), .Y(n1201) );
  AOI22X1TS U2069 ( .A0(n1196), .A1(readOutBus[548]), .B0(n1195), .B1(
        readOutBus[68]), .Y(n1200) );
  AOI22X1TS U2070 ( .A0(n1198), .A1(readOutBus[228]), .B0(n1197), .B1(
        readOutBus[388]), .Y(n1199) );
  NAND3XLTS U2071 ( .A(n1201), .B(n1200), .C(n1199), .Y(readOut[68]) );
  CLKBUFX2TS U2072 ( .A(n1238), .Y(n1212) );
  CLKBUFX2TS U2073 ( .A(n1239), .Y(n1211) );
  AOI22X1TS U2074 ( .A0(n1212), .A1(readOutBus[867]), .B0(n1211), .B1(
        readOutBus[707]), .Y(n1204) );
  CLKBUFX2TS U2075 ( .A(n1240), .Y(n1214) );
  CLKBUFX2TS U2076 ( .A(n1241), .Y(n1213) );
  AOI22X1TS U2077 ( .A0(n1214), .A1(readOutBus[547]), .B0(n1213), .B1(
        readOutBus[67]), .Y(n1203) );
  CLKBUFX2TS U2078 ( .A(n1242), .Y(n1216) );
  CLKBUFX2TS U2079 ( .A(n1243), .Y(n1215) );
  AOI22X1TS U2080 ( .A0(n1216), .A1(readOutBus[227]), .B0(n1215), .B1(
        readOutBus[387]), .Y(n1202) );
  NAND3XLTS U2081 ( .A(n1204), .B(n1203), .C(n1202), .Y(readOut[67]) );
  AOI22X1TS U2082 ( .A0(n1212), .A1(readOutBus[866]), .B0(n1211), .B1(
        readOutBus[706]), .Y(n1207) );
  AOI22X1TS U2083 ( .A0(n1214), .A1(readOutBus[546]), .B0(n1213), .B1(
        readOutBus[66]), .Y(n1206) );
  AOI22X1TS U2084 ( .A0(n1216), .A1(readOutBus[226]), .B0(n1215), .B1(
        readOutBus[386]), .Y(n1205) );
  NAND3XLTS U2085 ( .A(n1207), .B(n1206), .C(n1205), .Y(readOut[66]) );
  AOI22X1TS U2086 ( .A0(n1212), .A1(readOutBus[865]), .B0(n1211), .B1(
        readOutBus[705]), .Y(n1210) );
  AOI22X1TS U2087 ( .A0(n1214), .A1(readOutBus[545]), .B0(n1213), .B1(
        readOutBus[65]), .Y(n1209) );
  AOI22X1TS U2088 ( .A0(n1216), .A1(readOutBus[225]), .B0(n1215), .B1(
        readOutBus[385]), .Y(n1208) );
  NAND3XLTS U2089 ( .A(n1210), .B(n1209), .C(n1208), .Y(readOut[65]) );
  AOI22X1TS U2090 ( .A0(n1212), .A1(readOutBus[864]), .B0(n1211), .B1(
        readOutBus[704]), .Y(n1219) );
  AOI22X1TS U2091 ( .A0(n1214), .A1(readOutBus[544]), .B0(n1213), .B1(
        readOutBus[64]), .Y(n1218) );
  AOI22X1TS U2092 ( .A0(n1216), .A1(readOutBus[224]), .B0(n1215), .B1(
        readOutBus[384]), .Y(n1217) );
  NAND3XLTS U2093 ( .A(n1219), .B(n1218), .C(n1217), .Y(readOut[64]) );
  CLKBUFX2TS U2094 ( .A(n1238), .Y(n1230) );
  CLKBUFX2TS U2095 ( .A(n1239), .Y(n1229) );
  AOI22X1TS U2096 ( .A0(n1230), .A1(readOutBus[863]), .B0(n1229), .B1(
        readOutBus[703]), .Y(n1222) );
  CLKBUFX2TS U2097 ( .A(n1240), .Y(n1232) );
  CLKBUFX2TS U2098 ( .A(n1241), .Y(n1231) );
  AOI22X1TS U2099 ( .A0(n1232), .A1(readOutBus[543]), .B0(n1231), .B1(
        readOutBus[63]), .Y(n1221) );
  CLKBUFX2TS U2100 ( .A(n1242), .Y(n1234) );
  CLKBUFX2TS U2101 ( .A(n1243), .Y(n1233) );
  AOI22X1TS U2102 ( .A0(n1234), .A1(readOutBus[223]), .B0(n1233), .B1(
        readOutBus[383]), .Y(n1220) );
  NAND3XLTS U2103 ( .A(n1222), .B(n1221), .C(n1220), .Y(readOut[63]) );
  AOI22X1TS U2104 ( .A0(n1230), .A1(readOutBus[862]), .B0(n1229), .B1(
        readOutBus[702]), .Y(n1225) );
  AOI22X1TS U2105 ( .A0(n1232), .A1(readOutBus[542]), .B0(n1231), .B1(
        readOutBus[62]), .Y(n1224) );
  AOI22X1TS U2106 ( .A0(n1234), .A1(readOutBus[222]), .B0(n1233), .B1(
        readOutBus[382]), .Y(n1223) );
  NAND3XLTS U2107 ( .A(n1225), .B(n1224), .C(n1223), .Y(readOut[62]) );
  AOI22X1TS U2108 ( .A0(n1230), .A1(readOutBus[861]), .B0(n1229), .B1(
        readOutBus[701]), .Y(n1228) );
  AOI22X1TS U2109 ( .A0(n1232), .A1(readOutBus[541]), .B0(n1231), .B1(
        readOutBus[61]), .Y(n1227) );
  AOI22X1TS U2110 ( .A0(n1234), .A1(readOutBus[221]), .B0(n1233), .B1(
        readOutBus[381]), .Y(n1226) );
  NAND3XLTS U2111 ( .A(n1228), .B(n1227), .C(n1226), .Y(readOut[61]) );
  AOI22X1TS U2112 ( .A0(n1230), .A1(readOutBus[860]), .B0(n1229), .B1(
        readOutBus[700]), .Y(n1237) );
  AOI22X1TS U2113 ( .A0(n1232), .A1(readOutBus[540]), .B0(n1231), .B1(
        readOutBus[60]), .Y(n1236) );
  AOI22X1TS U2114 ( .A0(n1234), .A1(readOutBus[220]), .B0(n1233), .B1(
        readOutBus[380]), .Y(n1235) );
  NAND3XLTS U2115 ( .A(n1237), .B(n1236), .C(n1235), .Y(readOut[60]) );
  CLKBUFX2TS U2116 ( .A(n1238), .Y(n1254) );
  CLKBUFX2TS U2117 ( .A(n1239), .Y(n1253) );
  AOI22X1TS U2118 ( .A0(n1254), .A1(readOutBus[859]), .B0(n1253), .B1(
        readOutBus[699]), .Y(n1246) );
  CLKBUFX2TS U2119 ( .A(n1240), .Y(n1256) );
  CLKBUFX2TS U2120 ( .A(n1241), .Y(n1255) );
  AOI22X1TS U2121 ( .A0(n1256), .A1(readOutBus[539]), .B0(n1255), .B1(
        readOutBus[59]), .Y(n1245) );
  CLKBUFX2TS U2122 ( .A(n1242), .Y(n1258) );
  CLKBUFX2TS U2123 ( .A(n1243), .Y(n1257) );
  AOI22X1TS U2124 ( .A0(n1258), .A1(readOutBus[219]), .B0(n1257), .B1(
        readOutBus[379]), .Y(n1244) );
  NAND3XLTS U2125 ( .A(n1246), .B(n1245), .C(n1244), .Y(readOut[59]) );
  AOI22X1TS U2126 ( .A0(n1254), .A1(readOutBus[858]), .B0(n1253), .B1(
        readOutBus[698]), .Y(n1249) );
  AOI22X1TS U2127 ( .A0(n1256), .A1(readOutBus[538]), .B0(n1255), .B1(
        readOutBus[58]), .Y(n1248) );
  AOI22X1TS U2128 ( .A0(n1258), .A1(readOutBus[218]), .B0(n1257), .B1(
        readOutBus[378]), .Y(n1247) );
  NAND3XLTS U2129 ( .A(n1249), .B(n1248), .C(n1247), .Y(readOut[58]) );
  AOI22X1TS U2130 ( .A0(n1254), .A1(readOutBus[857]), .B0(n1253), .B1(
        readOutBus[697]), .Y(n1252) );
  AOI22X1TS U2131 ( .A0(n1256), .A1(readOutBus[537]), .B0(n1255), .B1(
        readOutBus[57]), .Y(n1251) );
  AOI22X1TS U2132 ( .A0(n1258), .A1(readOutBus[217]), .B0(n1257), .B1(
        readOutBus[377]), .Y(n1250) );
  NAND3XLTS U2133 ( .A(n1252), .B(n1251), .C(n1250), .Y(readOut[57]) );
  AOI22X1TS U2134 ( .A0(n1254), .A1(readOutBus[856]), .B0(n1253), .B1(
        readOutBus[696]), .Y(n1261) );
  AOI22X1TS U2135 ( .A0(n1256), .A1(readOutBus[536]), .B0(n1255), .B1(
        readOutBus[56]), .Y(n1260) );
  AOI22X1TS U2136 ( .A0(n1258), .A1(readOutBus[216]), .B0(n1257), .B1(
        readOutBus[376]), .Y(n1259) );
  NAND3XLTS U2137 ( .A(n1261), .B(n1260), .C(n1259), .Y(readOut[56]) );
  CLKBUFX2TS U2138 ( .A(n1298), .Y(n1272) );
  CLKBUFX2TS U2139 ( .A(n1299), .Y(n1271) );
  AOI22X1TS U2140 ( .A0(n1272), .A1(readOutBus[855]), .B0(n1271), .B1(
        readOutBus[695]), .Y(n1264) );
  CLKBUFX2TS U2141 ( .A(n1509), .Y(n1518) );
  CLKBUFX2TS U2142 ( .A(n1518), .Y(n1274) );
  CLKBUFX2TS U2143 ( .A(n1300), .Y(n1273) );
  AOI22X1TS U2144 ( .A0(n1274), .A1(readOutBus[535]), .B0(n1273), .B1(
        readOutBus[55]), .Y(n1263) );
  CLKBUFX2TS U2145 ( .A(n1511), .Y(n1520) );
  CLKBUFX2TS U2146 ( .A(n1520), .Y(n1276) );
  CLKBUFX2TS U2147 ( .A(n1301), .Y(n1275) );
  AOI22X1TS U2148 ( .A0(n1276), .A1(readOutBus[215]), .B0(n1275), .B1(
        readOutBus[375]), .Y(n1262) );
  NAND3XLTS U2149 ( .A(n1264), .B(n1263), .C(n1262), .Y(readOut[55]) );
  AOI22X1TS U2150 ( .A0(n1272), .A1(readOutBus[854]), .B0(n1271), .B1(
        readOutBus[694]), .Y(n1267) );
  AOI22X1TS U2151 ( .A0(n1274), .A1(readOutBus[534]), .B0(n1273), .B1(
        readOutBus[54]), .Y(n1266) );
  AOI22X1TS U2152 ( .A0(n1276), .A1(readOutBus[214]), .B0(n1275), .B1(
        readOutBus[374]), .Y(n1265) );
  NAND3XLTS U2153 ( .A(n1267), .B(n1266), .C(n1265), .Y(readOut[54]) );
  AOI22X1TS U2154 ( .A0(n1272), .A1(readOutBus[853]), .B0(n1271), .B1(
        readOutBus[693]), .Y(n1270) );
  AOI22X1TS U2155 ( .A0(n1274), .A1(readOutBus[533]), .B0(n1273), .B1(
        readOutBus[53]), .Y(n1269) );
  AOI22X1TS U2156 ( .A0(n1276), .A1(readOutBus[213]), .B0(n1275), .B1(
        readOutBus[373]), .Y(n1268) );
  NAND3XLTS U2157 ( .A(n1270), .B(n1269), .C(n1268), .Y(readOut[53]) );
  AOI22X1TS U2158 ( .A0(n1272), .A1(readOutBus[852]), .B0(n1271), .B1(
        readOutBus[692]), .Y(n1279) );
  AOI22X1TS U2159 ( .A0(n1274), .A1(readOutBus[532]), .B0(n1273), .B1(
        readOutBus[52]), .Y(n1278) );
  AOI22X1TS U2160 ( .A0(n1276), .A1(readOutBus[212]), .B0(n1275), .B1(
        readOutBus[372]), .Y(n1277) );
  NAND3XLTS U2161 ( .A(n1279), .B(n1278), .C(n1277), .Y(readOut[52]) );
  CLKBUFX2TS U2162 ( .A(n1298), .Y(n1290) );
  CLKBUFX2TS U2163 ( .A(n1299), .Y(n1289) );
  AOI22X1TS U2164 ( .A0(n1290), .A1(readOutBus[851]), .B0(n1289), .B1(
        readOutBus[691]), .Y(n1282) );
  CLKBUFX2TS U2165 ( .A(n1518), .Y(n1292) );
  CLKBUFX2TS U2166 ( .A(n1300), .Y(n1291) );
  AOI22X1TS U2167 ( .A0(n1292), .A1(readOutBus[531]), .B0(n1291), .B1(
        readOutBus[51]), .Y(n1281) );
  CLKBUFX2TS U2168 ( .A(n1520), .Y(n1294) );
  CLKBUFX2TS U2169 ( .A(n1301), .Y(n1293) );
  AOI22X1TS U2170 ( .A0(n1294), .A1(readOutBus[211]), .B0(n1293), .B1(
        readOutBus[371]), .Y(n1280) );
  NAND3XLTS U2171 ( .A(n1282), .B(n1281), .C(n1280), .Y(readOut[51]) );
  AOI22X1TS U2172 ( .A0(n1290), .A1(readOutBus[850]), .B0(n1289), .B1(
        readOutBus[690]), .Y(n1285) );
  AOI22X1TS U2173 ( .A0(n1292), .A1(readOutBus[530]), .B0(n1291), .B1(
        readOutBus[50]), .Y(n1284) );
  AOI22X1TS U2174 ( .A0(n1294), .A1(readOutBus[210]), .B0(n1293), .B1(
        readOutBus[370]), .Y(n1283) );
  NAND3XLTS U2175 ( .A(n1285), .B(n1284), .C(n1283), .Y(readOut[50]) );
  AOI22X1TS U2176 ( .A0(n1290), .A1(readOutBus[849]), .B0(n1289), .B1(
        readOutBus[689]), .Y(n1288) );
  AOI22X1TS U2177 ( .A0(n1292), .A1(readOutBus[529]), .B0(n1291), .B1(
        readOutBus[49]), .Y(n1287) );
  AOI22X1TS U2178 ( .A0(n1294), .A1(readOutBus[209]), .B0(n1293), .B1(
        readOutBus[369]), .Y(n1286) );
  NAND3XLTS U2179 ( .A(n1288), .B(n1287), .C(n1286), .Y(readOut[49]) );
  AOI22X1TS U2180 ( .A0(n1290), .A1(readOutBus[848]), .B0(n1289), .B1(
        readOutBus[688]), .Y(n1297) );
  AOI22X1TS U2181 ( .A0(n1292), .A1(readOutBus[528]), .B0(n1291), .B1(
        readOutBus[48]), .Y(n1296) );
  AOI22X1TS U2182 ( .A0(n1294), .A1(readOutBus[208]), .B0(n1293), .B1(
        readOutBus[368]), .Y(n1295) );
  NAND3XLTS U2183 ( .A(n1297), .B(n1296), .C(n1295), .Y(readOut[48]) );
  CLKBUFX2TS U2184 ( .A(n1298), .Y(n1312) );
  CLKBUFX2TS U2185 ( .A(n1299), .Y(n1311) );
  AOI22X1TS U2186 ( .A0(n1312), .A1(readOutBus[847]), .B0(n1311), .B1(
        readOutBus[687]), .Y(n1304) );
  CLKBUFX2TS U2187 ( .A(n1518), .Y(n1314) );
  CLKBUFX2TS U2188 ( .A(n1300), .Y(n1313) );
  AOI22X1TS U2189 ( .A0(n1314), .A1(readOutBus[527]), .B0(n1313), .B1(
        readOutBus[47]), .Y(n1303) );
  CLKBUFX2TS U2190 ( .A(n1520), .Y(n1316) );
  CLKBUFX2TS U2191 ( .A(n1301), .Y(n1315) );
  AOI22X1TS U2192 ( .A0(n1316), .A1(readOutBus[207]), .B0(n1315), .B1(
        readOutBus[367]), .Y(n1302) );
  NAND3XLTS U2193 ( .A(n1304), .B(n1303), .C(n1302), .Y(readOut[47]) );
  AOI22X1TS U2194 ( .A0(n1312), .A1(readOutBus[846]), .B0(n1311), .B1(
        readOutBus[686]), .Y(n1307) );
  AOI22X1TS U2195 ( .A0(n1314), .A1(readOutBus[526]), .B0(n1313), .B1(
        readOutBus[46]), .Y(n1306) );
  AOI22X1TS U2196 ( .A0(n1316), .A1(readOutBus[206]), .B0(n1315), .B1(
        readOutBus[366]), .Y(n1305) );
  NAND3XLTS U2197 ( .A(n1307), .B(n1306), .C(n1305), .Y(readOut[46]) );
  AOI22X1TS U2198 ( .A0(n1312), .A1(readOutBus[845]), .B0(n1311), .B1(
        readOutBus[685]), .Y(n1310) );
  AOI22X1TS U2199 ( .A0(n1314), .A1(readOutBus[525]), .B0(n1313), .B1(
        readOutBus[45]), .Y(n1309) );
  AOI22X1TS U2200 ( .A0(n1316), .A1(readOutBus[205]), .B0(n1315), .B1(
        readOutBus[365]), .Y(n1308) );
  NAND3XLTS U2201 ( .A(n1310), .B(n1309), .C(n1308), .Y(readOut[45]) );
  AOI22X1TS U2202 ( .A0(n1312), .A1(readOutBus[844]), .B0(n1311), .B1(
        readOutBus[684]), .Y(n1319) );
  AOI22X1TS U2203 ( .A0(n1314), .A1(readOutBus[524]), .B0(n1313), .B1(
        readOutBus[44]), .Y(n1318) );
  AOI22X1TS U2204 ( .A0(n1316), .A1(readOutBus[204]), .B0(n1315), .B1(
        readOutBus[364]), .Y(n1317) );
  NAND3XLTS U2205 ( .A(n1319), .B(n1318), .C(n1317), .Y(readOut[44]) );
  CLKBUFX2TS U2206 ( .A(n1356), .Y(n1330) );
  CLKBUFX2TS U2207 ( .A(n1357), .Y(n1329) );
  AOI22X1TS U2208 ( .A0(n1330), .A1(readOutBus[843]), .B0(n1329), .B1(
        readOutBus[683]), .Y(n1322) );
  CLKBUFX2TS U2209 ( .A(n1358), .Y(n1332) );
  CLKBUFX2TS U2210 ( .A(n1359), .Y(n1331) );
  AOI22X1TS U2211 ( .A0(n1332), .A1(readOutBus[523]), .B0(n1331), .B1(
        readOutBus[43]), .Y(n1321) );
  CLKBUFX2TS U2212 ( .A(n1360), .Y(n1334) );
  CLKBUFX2TS U2213 ( .A(n1361), .Y(n1333) );
  AOI22X1TS U2214 ( .A0(n1334), .A1(readOutBus[203]), .B0(n1333), .B1(
        readOutBus[363]), .Y(n1320) );
  NAND3XLTS U2215 ( .A(n1322), .B(n1321), .C(n1320), .Y(readOut[43]) );
  AOI22X1TS U2216 ( .A0(n1330), .A1(readOutBus[842]), .B0(n1329), .B1(
        readOutBus[682]), .Y(n1325) );
  AOI22X1TS U2217 ( .A0(n1332), .A1(readOutBus[522]), .B0(n1331), .B1(
        readOutBus[42]), .Y(n1324) );
  AOI22X1TS U2218 ( .A0(n1334), .A1(readOutBus[202]), .B0(n1333), .B1(
        readOutBus[362]), .Y(n1323) );
  NAND3XLTS U2219 ( .A(n1325), .B(n1324), .C(n1323), .Y(readOut[42]) );
  AOI22X1TS U2220 ( .A0(n1330), .A1(readOutBus[841]), .B0(n1329), .B1(
        readOutBus[681]), .Y(n1328) );
  AOI22X1TS U2221 ( .A0(n1332), .A1(readOutBus[521]), .B0(n1331), .B1(
        readOutBus[41]), .Y(n1327) );
  AOI22X1TS U2222 ( .A0(n1334), .A1(readOutBus[201]), .B0(n1333), .B1(
        readOutBus[361]), .Y(n1326) );
  NAND3XLTS U2223 ( .A(n1328), .B(n1327), .C(n1326), .Y(readOut[41]) );
  AOI22X1TS U2224 ( .A0(n1330), .A1(readOutBus[840]), .B0(n1329), .B1(
        readOutBus[680]), .Y(n1337) );
  AOI22X1TS U2225 ( .A0(n1332), .A1(readOutBus[520]), .B0(n1331), .B1(
        readOutBus[40]), .Y(n1336) );
  AOI22X1TS U2226 ( .A0(n1334), .A1(readOutBus[200]), .B0(n1333), .B1(
        readOutBus[360]), .Y(n1335) );
  NAND3XLTS U2227 ( .A(n1337), .B(n1336), .C(n1335), .Y(readOut[40]) );
  CLKBUFX2TS U2228 ( .A(n1356), .Y(n1348) );
  CLKBUFX2TS U2229 ( .A(n1357), .Y(n1347) );
  AOI22X1TS U2230 ( .A0(n1348), .A1(readOutBus[839]), .B0(n1347), .B1(
        readOutBus[679]), .Y(n1340) );
  CLKBUFX2TS U2231 ( .A(n1358), .Y(n1350) );
  CLKBUFX2TS U2232 ( .A(n1359), .Y(n1349) );
  AOI22X1TS U2233 ( .A0(n1350), .A1(readOutBus[519]), .B0(n1349), .B1(
        readOutBus[39]), .Y(n1339) );
  CLKBUFX2TS U2234 ( .A(n1360), .Y(n1352) );
  CLKBUFX2TS U2235 ( .A(n1361), .Y(n1351) );
  AOI22X1TS U2236 ( .A0(n1352), .A1(readOutBus[199]), .B0(n1351), .B1(
        readOutBus[359]), .Y(n1338) );
  NAND3XLTS U2237 ( .A(n1340), .B(n1339), .C(n1338), .Y(readOut[39]) );
  AOI22X1TS U2238 ( .A0(n1348), .A1(readOutBus[838]), .B0(n1347), .B1(
        readOutBus[678]), .Y(n1343) );
  AOI22X1TS U2239 ( .A0(n1350), .A1(readOutBus[518]), .B0(n1349), .B1(
        readOutBus[38]), .Y(n1342) );
  AOI22X1TS U2240 ( .A0(n1352), .A1(readOutBus[198]), .B0(n1351), .B1(
        readOutBus[358]), .Y(n1341) );
  NAND3XLTS U2241 ( .A(n1343), .B(n1342), .C(n1341), .Y(readOut[38]) );
  AOI22X1TS U2242 ( .A0(n1348), .A1(readOutBus[837]), .B0(n1347), .B1(
        readOutBus[677]), .Y(n1346) );
  AOI22X1TS U2243 ( .A0(n1350), .A1(readOutBus[517]), .B0(n1349), .B1(
        readOutBus[37]), .Y(n1345) );
  AOI22X1TS U2244 ( .A0(n1352), .A1(readOutBus[197]), .B0(n1351), .B1(
        readOutBus[357]), .Y(n1344) );
  NAND3XLTS U2245 ( .A(n1346), .B(n1345), .C(n1344), .Y(readOut[37]) );
  AOI22X1TS U2246 ( .A0(n1348), .A1(readOutBus[836]), .B0(n1347), .B1(
        readOutBus[676]), .Y(n1355) );
  AOI22X1TS U2247 ( .A0(n1350), .A1(readOutBus[516]), .B0(n1349), .B1(
        readOutBus[36]), .Y(n1354) );
  AOI22X1TS U2248 ( .A0(n1352), .A1(readOutBus[196]), .B0(n1351), .B1(
        readOutBus[356]), .Y(n1353) );
  NAND3XLTS U2249 ( .A(n1355), .B(n1354), .C(n1353), .Y(readOut[36]) );
  CLKBUFX2TS U2250 ( .A(n1356), .Y(n1372) );
  CLKBUFX2TS U2251 ( .A(n1357), .Y(n1371) );
  AOI22X1TS U2252 ( .A0(n1372), .A1(readOutBus[835]), .B0(n1371), .B1(
        readOutBus[675]), .Y(n1364) );
  CLKBUFX2TS U2253 ( .A(n1358), .Y(n1374) );
  CLKBUFX2TS U2254 ( .A(n1359), .Y(n1373) );
  AOI22X1TS U2255 ( .A0(n1374), .A1(readOutBus[515]), .B0(n1373), .B1(
        readOutBus[35]), .Y(n1363) );
  CLKBUFX2TS U2256 ( .A(n1360), .Y(n1376) );
  CLKBUFX2TS U2257 ( .A(n1361), .Y(n1375) );
  AOI22X1TS U2258 ( .A0(n1376), .A1(readOutBus[195]), .B0(n1375), .B1(
        readOutBus[355]), .Y(n1362) );
  NAND3XLTS U2259 ( .A(n1364), .B(n1363), .C(n1362), .Y(readOut[35]) );
  AOI22X1TS U2260 ( .A0(n1372), .A1(readOutBus[834]), .B0(n1371), .B1(
        readOutBus[674]), .Y(n1367) );
  AOI22X1TS U2261 ( .A0(n1374), .A1(readOutBus[514]), .B0(n1373), .B1(
        readOutBus[34]), .Y(n1366) );
  AOI22X1TS U2262 ( .A0(n1376), .A1(readOutBus[194]), .B0(n1375), .B1(
        readOutBus[354]), .Y(n1365) );
  NAND3XLTS U2263 ( .A(n1367), .B(n1366), .C(n1365), .Y(readOut[34]) );
  AOI22X1TS U2264 ( .A0(n1372), .A1(readOutBus[833]), .B0(n1371), .B1(
        readOutBus[673]), .Y(n1370) );
  AOI22X1TS U2265 ( .A0(n1374), .A1(readOutBus[513]), .B0(n1373), .B1(
        readOutBus[33]), .Y(n1369) );
  AOI22X1TS U2266 ( .A0(n1376), .A1(readOutBus[193]), .B0(n1375), .B1(
        readOutBus[353]), .Y(n1368) );
  NAND3XLTS U2267 ( .A(n1370), .B(n1369), .C(n1368), .Y(readOut[33]) );
  AOI22X1TS U2268 ( .A0(n1372), .A1(readOutBus[832]), .B0(n1371), .B1(
        readOutBus[672]), .Y(n1379) );
  AOI22X1TS U2269 ( .A0(n1374), .A1(readOutBus[512]), .B0(n1373), .B1(
        readOutBus[32]), .Y(n1378) );
  AOI22X1TS U2270 ( .A0(n1376), .A1(readOutBus[192]), .B0(n1375), .B1(
        readOutBus[352]), .Y(n1377) );
  NAND3XLTS U2271 ( .A(n1379), .B(n1378), .C(n1377), .Y(readOut[32]) );
  CLKBUFX2TS U2272 ( .A(n1416), .Y(n1390) );
  CLKBUFX2TS U2273 ( .A(n1417), .Y(n1389) );
  AOI22X1TS U2274 ( .A0(n1390), .A1(readOutBus[831]), .B0(n1389), .B1(
        readOutBus[671]), .Y(n1382) );
  CLKBUFX2TS U2275 ( .A(n1418), .Y(n1392) );
  CLKBUFX2TS U2276 ( .A(n1419), .Y(n1391) );
  AOI22X1TS U2277 ( .A0(n1392), .A1(readOutBus[511]), .B0(n1391), .B1(
        readOutBus[31]), .Y(n1381) );
  CLKBUFX2TS U2278 ( .A(n1420), .Y(n1394) );
  CLKBUFX2TS U2279 ( .A(n1421), .Y(n1393) );
  AOI22X1TS U2280 ( .A0(n1394), .A1(readOutBus[191]), .B0(n1393), .B1(
        readOutBus[351]), .Y(n1380) );
  NAND3XLTS U2281 ( .A(n1382), .B(n1381), .C(n1380), .Y(readOut[31]) );
  AOI22X1TS U2282 ( .A0(n1390), .A1(readOutBus[830]), .B0(n1389), .B1(
        readOutBus[670]), .Y(n1385) );
  AOI22X1TS U2283 ( .A0(n1392), .A1(readOutBus[510]), .B0(n1391), .B1(
        readOutBus[30]), .Y(n1384) );
  AOI22X1TS U2284 ( .A0(n1394), .A1(readOutBus[190]), .B0(n1393), .B1(
        readOutBus[350]), .Y(n1383) );
  NAND3XLTS U2285 ( .A(n1385), .B(n1384), .C(n1383), .Y(readOut[30]) );
  AOI22X1TS U2286 ( .A0(n1390), .A1(readOutBus[829]), .B0(n1389), .B1(
        readOutBus[669]), .Y(n1388) );
  AOI22X1TS U2287 ( .A0(n1392), .A1(readOutBus[509]), .B0(n1391), .B1(
        readOutBus[29]), .Y(n1387) );
  AOI22X1TS U2288 ( .A0(n1394), .A1(readOutBus[189]), .B0(n1393), .B1(
        readOutBus[349]), .Y(n1386) );
  NAND3XLTS U2289 ( .A(n1388), .B(n1387), .C(n1386), .Y(readOut[29]) );
  AOI22X1TS U2290 ( .A0(n1390), .A1(readOutBus[828]), .B0(n1389), .B1(
        readOutBus[668]), .Y(n1397) );
  AOI22X1TS U2291 ( .A0(n1392), .A1(readOutBus[508]), .B0(n1391), .B1(
        readOutBus[28]), .Y(n1396) );
  AOI22X1TS U2292 ( .A0(n1394), .A1(readOutBus[188]), .B0(n1393), .B1(
        readOutBus[348]), .Y(n1395) );
  NAND3XLTS U2293 ( .A(n1397), .B(n1396), .C(n1395), .Y(readOut[28]) );
  CLKBUFX2TS U2294 ( .A(n1416), .Y(n1408) );
  CLKBUFX2TS U2295 ( .A(n1417), .Y(n1407) );
  AOI22X1TS U2296 ( .A0(n1408), .A1(readOutBus[827]), .B0(n1407), .B1(
        readOutBus[667]), .Y(n1400) );
  CLKBUFX2TS U2297 ( .A(n1418), .Y(n1410) );
  CLKBUFX2TS U2298 ( .A(n1419), .Y(n1409) );
  AOI22X1TS U2299 ( .A0(n1410), .A1(readOutBus[507]), .B0(n1409), .B1(
        readOutBus[27]), .Y(n1399) );
  CLKBUFX2TS U2300 ( .A(n1420), .Y(n1412) );
  CLKBUFX2TS U2301 ( .A(n1421), .Y(n1411) );
  AOI22X1TS U2302 ( .A0(n1412), .A1(readOutBus[187]), .B0(n1411), .B1(
        readOutBus[347]), .Y(n1398) );
  NAND3XLTS U2303 ( .A(n1400), .B(n1399), .C(n1398), .Y(readOut[27]) );
  AOI22X1TS U2304 ( .A0(n1408), .A1(readOutBus[826]), .B0(n1407), .B1(
        readOutBus[666]), .Y(n1403) );
  AOI22X1TS U2305 ( .A0(n1410), .A1(readOutBus[506]), .B0(n1409), .B1(
        readOutBus[26]), .Y(n1402) );
  AOI22X1TS U2306 ( .A0(n1412), .A1(readOutBus[186]), .B0(n1411), .B1(
        readOutBus[346]), .Y(n1401) );
  NAND3XLTS U2307 ( .A(n1403), .B(n1402), .C(n1401), .Y(readOut[26]) );
  AOI22X1TS U2308 ( .A0(n1408), .A1(readOutBus[825]), .B0(n1407), .B1(
        readOutBus[665]), .Y(n1406) );
  AOI22X1TS U2309 ( .A0(n1410), .A1(readOutBus[505]), .B0(n1409), .B1(
        readOutBus[25]), .Y(n1405) );
  AOI22X1TS U2310 ( .A0(n1412), .A1(readOutBus[185]), .B0(n1411), .B1(
        readOutBus[345]), .Y(n1404) );
  NAND3XLTS U2311 ( .A(n1406), .B(n1405), .C(n1404), .Y(readOut[25]) );
  AOI22X1TS U2312 ( .A0(n1408), .A1(readOutBus[824]), .B0(n1407), .B1(
        readOutBus[664]), .Y(n1415) );
  AOI22X1TS U2313 ( .A0(n1410), .A1(readOutBus[504]), .B0(n1409), .B1(
        readOutBus[24]), .Y(n1414) );
  AOI22X1TS U2314 ( .A0(n1412), .A1(readOutBus[184]), .B0(n1411), .B1(
        readOutBus[344]), .Y(n1413) );
  NAND3XLTS U2315 ( .A(n1415), .B(n1414), .C(n1413), .Y(readOut[24]) );
  CLKBUFX2TS U2316 ( .A(n1416), .Y(n1432) );
  CLKBUFX2TS U2317 ( .A(n1417), .Y(n1431) );
  AOI22X1TS U2318 ( .A0(n1432), .A1(readOutBus[823]), .B0(n1431), .B1(
        readOutBus[663]), .Y(n1424) );
  CLKBUFX2TS U2319 ( .A(n1418), .Y(n1434) );
  CLKBUFX2TS U2320 ( .A(n1419), .Y(n1433) );
  AOI22X1TS U2321 ( .A0(n1434), .A1(readOutBus[503]), .B0(n1433), .B1(
        readOutBus[23]), .Y(n1423) );
  CLKBUFX2TS U2322 ( .A(n1420), .Y(n1436) );
  CLKBUFX2TS U2323 ( .A(n1421), .Y(n1435) );
  AOI22X1TS U2324 ( .A0(n1436), .A1(readOutBus[183]), .B0(n1435), .B1(
        readOutBus[343]), .Y(n1422) );
  NAND3XLTS U2325 ( .A(n1424), .B(n1423), .C(n1422), .Y(readOut[23]) );
  AOI22X1TS U2326 ( .A0(n1432), .A1(readOutBus[822]), .B0(n1431), .B1(
        readOutBus[662]), .Y(n1427) );
  AOI22X1TS U2327 ( .A0(n1434), .A1(readOutBus[502]), .B0(n1433), .B1(
        readOutBus[22]), .Y(n1426) );
  AOI22X1TS U2328 ( .A0(n1436), .A1(readOutBus[182]), .B0(n1435), .B1(
        readOutBus[342]), .Y(n1425) );
  NAND3XLTS U2329 ( .A(n1427), .B(n1426), .C(n1425), .Y(readOut[22]) );
  AOI22X1TS U2330 ( .A0(n1432), .A1(readOutBus[821]), .B0(n1431), .B1(
        readOutBus[661]), .Y(n1430) );
  AOI22X1TS U2331 ( .A0(n1434), .A1(readOutBus[501]), .B0(n1433), .B1(
        readOutBus[21]), .Y(n1429) );
  AOI22X1TS U2332 ( .A0(n1436), .A1(readOutBus[181]), .B0(n1435), .B1(
        readOutBus[341]), .Y(n1428) );
  NAND3XLTS U2333 ( .A(n1430), .B(n1429), .C(n1428), .Y(readOut[21]) );
  AOI22X1TS U2334 ( .A0(n1432), .A1(readOutBus[820]), .B0(n1431), .B1(
        readOutBus[660]), .Y(n1439) );
  AOI22X1TS U2335 ( .A0(n1434), .A1(readOutBus[500]), .B0(n1433), .B1(
        readOutBus[20]), .Y(n1438) );
  AOI22X1TS U2336 ( .A0(n1436), .A1(readOutBus[180]), .B0(n1435), .B1(
        readOutBus[340]), .Y(n1437) );
  NAND3XLTS U2337 ( .A(n1439), .B(n1438), .C(n1437), .Y(readOut[20]) );
  CLKBUFX2TS U2338 ( .A(n1476), .Y(n1450) );
  CLKBUFX2TS U2339 ( .A(n1477), .Y(n1449) );
  AOI22X1TS U2340 ( .A0(n1450), .A1(readOutBus[819]), .B0(n1449), .B1(
        readOutBus[659]), .Y(n1442) );
  CLKBUFX2TS U2341 ( .A(n1478), .Y(n1452) );
  CLKBUFX2TS U2342 ( .A(n1479), .Y(n1451) );
  AOI22X1TS U2343 ( .A0(n1452), .A1(readOutBus[499]), .B0(n1451), .B1(
        readOutBus[19]), .Y(n1441) );
  CLKBUFX2TS U2344 ( .A(n1480), .Y(n1454) );
  CLKBUFX2TS U2345 ( .A(n1481), .Y(n1453) );
  AOI22X1TS U2346 ( .A0(n1454), .A1(readOutBus[179]), .B0(n1453), .B1(
        readOutBus[339]), .Y(n1440) );
  NAND3XLTS U2347 ( .A(n1442), .B(n1441), .C(n1440), .Y(readOut[19]) );
  AOI22X1TS U2348 ( .A0(n1450), .A1(readOutBus[818]), .B0(n1449), .B1(
        readOutBus[658]), .Y(n1445) );
  AOI22X1TS U2349 ( .A0(n1452), .A1(readOutBus[498]), .B0(n1451), .B1(
        readOutBus[18]), .Y(n1444) );
  AOI22X1TS U2350 ( .A0(n1454), .A1(readOutBus[178]), .B0(n1453), .B1(
        readOutBus[338]), .Y(n1443) );
  NAND3XLTS U2351 ( .A(n1445), .B(n1444), .C(n1443), .Y(readOut[18]) );
  AOI22X1TS U2352 ( .A0(n1450), .A1(readOutBus[817]), .B0(n1449), .B1(
        readOutBus[657]), .Y(n1448) );
  AOI22X1TS U2353 ( .A0(n1452), .A1(readOutBus[497]), .B0(n1451), .B1(
        readOutBus[17]), .Y(n1447) );
  AOI22X1TS U2354 ( .A0(n1454), .A1(readOutBus[177]), .B0(n1453), .B1(
        readOutBus[337]), .Y(n1446) );
  NAND3XLTS U2355 ( .A(n1448), .B(n1447), .C(n1446), .Y(readOut[17]) );
  AOI22X1TS U2356 ( .A0(n1450), .A1(readOutBus[816]), .B0(n1449), .B1(
        readOutBus[656]), .Y(n1457) );
  AOI22X1TS U2357 ( .A0(n1452), .A1(readOutBus[496]), .B0(n1451), .B1(
        readOutBus[16]), .Y(n1456) );
  AOI22X1TS U2358 ( .A0(n1454), .A1(readOutBus[176]), .B0(n1453), .B1(
        readOutBus[336]), .Y(n1455) );
  NAND3XLTS U2359 ( .A(n1457), .B(n1456), .C(n1455), .Y(readOut[16]) );
  CLKBUFX2TS U2360 ( .A(n1476), .Y(n1468) );
  CLKBUFX2TS U2361 ( .A(n1477), .Y(n1467) );
  AOI22X1TS U2362 ( .A0(n1468), .A1(readOutBus[815]), .B0(n1467), .B1(
        readOutBus[655]), .Y(n1460) );
  CLKBUFX2TS U2363 ( .A(n1478), .Y(n1470) );
  CLKBUFX2TS U2364 ( .A(n1479), .Y(n1469) );
  AOI22X1TS U2365 ( .A0(n1470), .A1(readOutBus[495]), .B0(n1469), .B1(
        readOutBus[15]), .Y(n1459) );
  CLKBUFX2TS U2366 ( .A(n1480), .Y(n1472) );
  CLKBUFX2TS U2367 ( .A(n1481), .Y(n1471) );
  AOI22X1TS U2368 ( .A0(n1472), .A1(readOutBus[175]), .B0(n1471), .B1(
        readOutBus[335]), .Y(n1458) );
  NAND3XLTS U2369 ( .A(n1460), .B(n1459), .C(n1458), .Y(readOut[15]) );
  AOI22X1TS U2370 ( .A0(n1468), .A1(readOutBus[814]), .B0(n1467), .B1(
        readOutBus[654]), .Y(n1463) );
  AOI22X1TS U2371 ( .A0(n1470), .A1(readOutBus[494]), .B0(n1469), .B1(
        readOutBus[14]), .Y(n1462) );
  AOI22X1TS U2372 ( .A0(n1472), .A1(readOutBus[174]), .B0(n1471), .B1(
        readOutBus[334]), .Y(n1461) );
  NAND3XLTS U2373 ( .A(n1463), .B(n1462), .C(n1461), .Y(readOut[14]) );
  AOI22X1TS U2374 ( .A0(n1468), .A1(readOutBus[813]), .B0(n1467), .B1(
        readOutBus[653]), .Y(n1466) );
  AOI22X1TS U2375 ( .A0(n1470), .A1(readOutBus[493]), .B0(n1469), .B1(
        readOutBus[13]), .Y(n1465) );
  AOI22X1TS U2376 ( .A0(n1472), .A1(readOutBus[173]), .B0(n1471), .B1(
        readOutBus[333]), .Y(n1464) );
  NAND3XLTS U2377 ( .A(n1466), .B(n1465), .C(n1464), .Y(readOut[13]) );
  AOI22X1TS U2378 ( .A0(n1468), .A1(readOutBus[812]), .B0(n1467), .B1(
        readOutBus[652]), .Y(n1475) );
  AOI22X1TS U2379 ( .A0(n1470), .A1(readOutBus[492]), .B0(n1469), .B1(
        readOutBus[12]), .Y(n1474) );
  AOI22X1TS U2380 ( .A0(n1472), .A1(readOutBus[172]), .B0(n1471), .B1(
        readOutBus[332]), .Y(n1473) );
  NAND3XLTS U2381 ( .A(n1475), .B(n1474), .C(n1473), .Y(readOut[12]) );
  CLKBUFX2TS U2382 ( .A(n1476), .Y(n1492) );
  CLKBUFX2TS U2383 ( .A(n1477), .Y(n1491) );
  AOI22X1TS U2384 ( .A0(n1492), .A1(readOutBus[811]), .B0(n1491), .B1(
        readOutBus[651]), .Y(n1484) );
  CLKBUFX2TS U2385 ( .A(n1478), .Y(n1494) );
  CLKBUFX2TS U2386 ( .A(n1479), .Y(n1493) );
  AOI22X1TS U2387 ( .A0(n1494), .A1(readOutBus[491]), .B0(n1493), .B1(
        readOutBus[11]), .Y(n1483) );
  CLKBUFX2TS U2388 ( .A(n1480), .Y(n1496) );
  CLKBUFX2TS U2389 ( .A(n1481), .Y(n1495) );
  AOI22X1TS U2390 ( .A0(n1496), .A1(readOutBus[171]), .B0(n1495), .B1(
        readOutBus[331]), .Y(n1482) );
  NAND3XLTS U2391 ( .A(n1484), .B(n1483), .C(n1482), .Y(readOut[11]) );
  AOI22X1TS U2392 ( .A0(n1492), .A1(readOutBus[810]), .B0(n1491), .B1(
        readOutBus[650]), .Y(n1487) );
  AOI22X1TS U2393 ( .A0(n1494), .A1(readOutBus[490]), .B0(n1493), .B1(
        readOutBus[10]), .Y(n1486) );
  AOI22X1TS U2394 ( .A0(n1496), .A1(readOutBus[170]), .B0(n1495), .B1(
        readOutBus[330]), .Y(n1485) );
  NAND3XLTS U2395 ( .A(n1487), .B(n1486), .C(n1485), .Y(readOut[10]) );
  AOI22X1TS U2396 ( .A0(n1492), .A1(readOutBus[809]), .B0(n1491), .B1(
        readOutBus[649]), .Y(n1490) );
  AOI22X1TS U2397 ( .A0(n1494), .A1(readOutBus[489]), .B0(n1493), .B1(
        readOutBus[9]), .Y(n1489) );
  AOI22X1TS U2398 ( .A0(n1496), .A1(readOutBus[169]), .B0(n1495), .B1(
        readOutBus[329]), .Y(n1488) );
  NAND3XLTS U2399 ( .A(n1490), .B(n1489), .C(n1488), .Y(readOut[9]) );
  AOI22X1TS U2400 ( .A0(n1492), .A1(readOutBus[808]), .B0(n1491), .B1(
        readOutBus[648]), .Y(n1499) );
  AOI22X1TS U2401 ( .A0(n1494), .A1(readOutBus[488]), .B0(n1493), .B1(
        readOutBus[8]), .Y(n1498) );
  AOI22X1TS U2402 ( .A0(n1496), .A1(readOutBus[168]), .B0(n1495), .B1(
        readOutBus[328]), .Y(n1497) );
  NAND3XLTS U2403 ( .A(n1499), .B(n1498), .C(n1497), .Y(readOut[8]) );
  AOI22X1TS U2404 ( .A0(n1540), .A1(readOutBus[807]), .B0(n1539), .B1(
        readOutBus[647]), .Y(n1502) );
  AOI22X1TS U2405 ( .A0(n1542), .A1(readOutBus[487]), .B0(n1541), .B1(
        readOutBus[7]), .Y(n1501) );
  AOI22X1TS U2406 ( .A0(n1544), .A1(readOutBus[167]), .B0(n1543), .B1(
        readOutBus[327]), .Y(n1500) );
  NAND3XLTS U2407 ( .A(n1502), .B(n1501), .C(n1500), .Y(readOut[7]) );
  AOI22X1TS U2408 ( .A0(n1540), .A1(readOutBus[806]), .B0(n1539), .B1(
        readOutBus[646]), .Y(n1505) );
  AOI22X1TS U2409 ( .A0(n1542), .A1(readOutBus[486]), .B0(n1541), .B1(
        readOutBus[6]), .Y(n1504) );
  AOI22X1TS U2410 ( .A0(n1544), .A1(readOutBus[166]), .B0(n1543), .B1(
        readOutBus[326]), .Y(n1503) );
  NAND3XLTS U2411 ( .A(n1505), .B(n1504), .C(n1503), .Y(readOut[6]) );
  AOI22X1TS U2412 ( .A0(n1507), .A1(readOutBus[805]), .B0(n1506), .B1(
        readOutBus[645]), .Y(n1514) );
  AOI22X1TS U2413 ( .A0(n1509), .A1(readOutBus[485]), .B0(n1508), .B1(
        readOutBus[5]), .Y(n1513) );
  AOI22X1TS U2414 ( .A0(n1511), .A1(readOutBus[165]), .B0(n1510), .B1(
        readOutBus[325]), .Y(n1512) );
  NAND3XLTS U2415 ( .A(n1514), .B(n1513), .C(n1512), .Y(readOut[5]) );
  AOI22X1TS U2416 ( .A0(n1516), .A1(readOutBus[804]), .B0(n1515), .B1(
        readOutBus[644]), .Y(n1523) );
  AOI22X1TS U2417 ( .A0(n1518), .A1(readOutBus[484]), .B0(n1517), .B1(
        readOutBus[4]), .Y(n1522) );
  AOI22X1TS U2418 ( .A0(n1520), .A1(readOutBus[164]), .B0(n1519), .B1(
        readOutBus[324]), .Y(n1521) );
  NAND3XLTS U2419 ( .A(n1523), .B(n1522), .C(n1521), .Y(readOut[4]) );
  AOI22X1TS U2420 ( .A0(n1531), .A1(readOutBus[803]), .B0(n1530), .B1(
        readOutBus[643]), .Y(n1526) );
  AOI22X1TS U2421 ( .A0(n1533), .A1(readOutBus[483]), .B0(n1532), .B1(
        readOutBus[3]), .Y(n1525) );
  AOI22X1TS U2422 ( .A0(n1535), .A1(readOutBus[163]), .B0(n1534), .B1(
        readOutBus[323]), .Y(n1524) );
  NAND3XLTS U2423 ( .A(n1526), .B(n1525), .C(n1524), .Y(readOut[3]) );
  AOI22X1TS U2424 ( .A0(n1531), .A1(readOutBus[802]), .B0(n1530), .B1(
        readOutBus[642]), .Y(n1529) );
  AOI22X1TS U2425 ( .A0(n1533), .A1(readOutBus[482]), .B0(n1532), .B1(
        readOutBus[2]), .Y(n1528) );
  AOI22X1TS U2426 ( .A0(n1535), .A1(readOutBus[162]), .B0(n1534), .B1(
        readOutBus[322]), .Y(n1527) );
  NAND3XLTS U2427 ( .A(n1529), .B(n1528), .C(n1527), .Y(readOut[2]) );
  AOI22X1TS U2428 ( .A0(n1531), .A1(readOutBus[801]), .B0(n1530), .B1(
        readOutBus[641]), .Y(n1538) );
  AOI22X1TS U2429 ( .A0(n1533), .A1(readOutBus[481]), .B0(n1532), .B1(
        readOutBus[1]), .Y(n1537) );
  AOI22X1TS U2430 ( .A0(n1535), .A1(readOutBus[161]), .B0(n1534), .B1(
        readOutBus[321]), .Y(n1536) );
  NAND3XLTS U2431 ( .A(n1538), .B(n1537), .C(n1536), .Y(readOut[1]) );
  AOI22X1TS U2432 ( .A0(n1540), .A1(readOutBus[800]), .B0(n1539), .B1(
        readOutBus[640]), .Y(n1547) );
  AOI22X1TS U2433 ( .A0(n1542), .A1(readOutBus[480]), .B0(n1541), .B1(
        readOutBus[0]), .Y(n1546) );
  AOI22X1TS U2434 ( .A0(n1544), .A1(readOutBus[160]), .B0(n1543), .B1(
        readOutBus[320]), .Y(n1545) );
  NAND3XLTS U2435 ( .A(n1547), .B(n1546), .C(n1545), .Y(readOut[0]) );
endmodule

