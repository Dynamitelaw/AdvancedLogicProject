
module InputQueueRegister ( clk, resetInputQueue, resetBuffer, pixelValue, 
        dequeue, writeBufferEnable, finished, indexOut, queueEmpty );
  output [9:0] indexOut;
  input clk, resetInputQueue, resetBuffer, pixelValue, dequeue,
         writeBufferEnable;
  output finished, queueEmpty;
  wire   N89, N90, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N126, N127, n85, n86, n87, n88, n890, n900, n91, n92, n93, n94, n95,
         n96, n97, n980, n990, n1000, n1010, n1020, n1030, n1040, n1050, n1060,
         n1070, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n1260, n1270, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n178, n181, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553;
  wire   [9:0] queueEndPointerBuffer;
  wire   [9:0] queueEndPointer;
  wire   [69:0] queueRegister;
  wire   [69:0] queueRegisterBuffer;
  wire   [9:0] indexCounter;
  wire   [9:0] queueFrontPointerBuffer;

  DFFRX4TS queueEndPointer_reg_2_ ( .D(n181), .CK(clk), .RN(n553), .Q(n478), 
        .QN(n499) );
  DFFNSRX1TS indexCounter_reg_6_ ( .D(n980), .CKN(clk), .SN(1'b1), .RN(n484), 
        .Q(indexCounter[6]), .QN(n493) );
  DFFNSRX1TS indexCounter_reg_7_ ( .D(n97), .CKN(clk), .SN(1'b1), .RN(n480), 
        .Q(indexCounter[7]), .QN(n534) );
  DFFNSRX1TS indexCounter_reg_8_ ( .D(n96), .CKN(clk), .SN(1'b1), .RN(n553), 
        .Q(indexCounter[8]), .QN(n533) );
  DFFNSRX1TS indexCounter_reg_5_ ( .D(n990), .CKN(clk), .SN(1'b1), .RN(n220), 
        .Q(indexCounter[5]), .QN(n532) );
  DFFNSRX1TS indexCounter_reg_2_ ( .D(n1020), .CKN(clk), .SN(1'b1), .RN(n219), 
        .Q(indexCounter[2]), .QN(n531) );
  DFFNSRX1TS indexCounter_reg_3_ ( .D(n1010), .CKN(clk), .SN(1'b1), .RN(n480), 
        .Q(indexCounter[3]), .QN(n529) );
  DFFNSRX1TS indexCounter_reg_0_ ( .D(n1040), .CKN(clk), .SN(1'b1), .RN(n479), 
        .Q(indexCounter[0]), .QN(n530) );
  DFFNSRX1TS indexCounter_reg_4_ ( .D(n1000), .CKN(clk), .SN(1'b1), .RN(n484), 
        .Q(indexCounter[4]), .QN(n495) );
  DFFNSRX1TS indexCounter_reg_1_ ( .D(n1030), .CKN(clk), .SN(1'b1), .RN(n480), 
        .Q(indexCounter[1]), .QN(n494) );
  DFFSX4TS queueEndPointer_reg_1_ ( .D(n497), .CK(clk), .SN(n553), .Q(n526), 
        .QN(queueEndPointer[1]) );
  DFFSX4TS queueEndPointer_reg_8_ ( .D(n511), .CK(clk), .SN(n479), .Q(n527), 
        .QN(queueEndPointer[8]) );
  DFFSX4TS queueEndPointer_reg_7_ ( .D(n510), .CK(clk), .SN(n479), .Q(n522), 
        .QN(queueEndPointer[7]) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_5_ ( .D(n890), .CKN(n488), .SN(1'b1), 
        .RN(n482), .Q(queueFrontPointerBuffer[5]), .QN(n507) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_8_ ( .D(n86), .CKN(n486), .SN(1'b1), 
        .RN(n483), .Q(queueFrontPointerBuffer[8]), .QN(n506) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_7_ ( .D(n87), .CKN(n477), .SN(1'b1), 
        .RN(n482), .Q(queueFrontPointerBuffer[7]), .QN(n505) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_9_ ( .D(n85), .CKN(n486), .SN(1'b1), 
        .RN(n483), .Q(queueFrontPointerBuffer[9]), .QN(n504) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_3_ ( .D(n91), .CKN(n488), .SN(1'b1), 
        .RN(n482), .Q(queueFrontPointerBuffer[3]), .QN(n503) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_6_ ( .D(n88), .CKN(n477), .SN(1'b1), 
        .RN(n483), .QN(n502) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_4_ ( .D(n900), .CKN(n487), .SN(1'b1), 
        .RN(n481), .QN(n501) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_2_ ( .D(n92), .CKN(n485), .SN(1'b1), 
        .RN(n481), .Q(queueFrontPointerBuffer[2]), .QN(n500) );
  DFFQX1TS queueRegisterBuffer_reg_5__6_ ( .D(queueRegister[56]), .CK(n544), 
        .Q(queueRegisterBuffer[56]) );
  DFFQX1TS queueRegisterBuffer_reg_5__7_ ( .D(queueRegister[57]), .CK(n544), 
        .Q(queueRegisterBuffer[57]) );
  DFFQX1TS queueRegisterBuffer_reg_5__8_ ( .D(queueRegister[58]), .CK(n544), 
        .Q(queueRegisterBuffer[58]) );
  DFFQX1TS queueRegisterBuffer_reg_4__9_ ( .D(queueRegister[49]), .CK(n549), 
        .Q(queueRegisterBuffer[49]) );
  DFFQX1TS queueRegisterBuffer_reg_5__9_ ( .D(queueRegister[59]), .CK(n542), 
        .Q(queueRegisterBuffer[59]) );
  DFFQX1TS queueRegisterBuffer_reg_5__0_ ( .D(queueRegister[50]), .CK(n542), 
        .Q(queueRegisterBuffer[50]) );
  DFFQX1TS queueRegisterBuffer_reg_5__1_ ( .D(queueRegister[51]), .CK(n542), 
        .Q(queueRegisterBuffer[51]) );
  DFFQX1TS queueRegisterBuffer_reg_5__2_ ( .D(queueRegister[52]), .CK(n543), 
        .Q(queueRegisterBuffer[52]) );
  DFFQX1TS queueRegisterBuffer_reg_5__3_ ( .D(queueRegister[53]), .CK(n543), 
        .Q(queueRegisterBuffer[53]) );
  DFFQX1TS queueRegisterBuffer_reg_5__4_ ( .D(queueRegister[54]), .CK(n543), 
        .Q(queueRegisterBuffer[54]) );
  DFFQX1TS queueRegisterBuffer_reg_5__5_ ( .D(queueRegister[55]), .CK(n543), 
        .Q(queueRegisterBuffer[55]) );
  DFFQX1TS queueRegisterBuffer_reg_4__0_ ( .D(queueRegister[40]), .CK(n550), 
        .Q(queueRegisterBuffer[40]) );
  DFFQX1TS queueRegisterBuffer_reg_4__1_ ( .D(queueRegister[41]), .CK(n550), 
        .Q(queueRegisterBuffer[41]) );
  DFFQX1TS queueRegisterBuffer_reg_4__2_ ( .D(queueRegister[42]), .CK(n550), 
        .Q(queueRegisterBuffer[42]) );
  DFFQX1TS queueRegisterBuffer_reg_4__3_ ( .D(queueRegister[43]), .CK(n550), 
        .Q(queueRegisterBuffer[43]) );
  DFFQX1TS queueRegisterBuffer_reg_4__4_ ( .D(queueRegister[44]), .CK(n551), 
        .Q(queueRegisterBuffer[44]) );
  DFFQX1TS queueRegisterBuffer_reg_4__5_ ( .D(queueRegister[45]), .CK(n551), 
        .Q(queueRegisterBuffer[45]) );
  DFFQX1TS queueRegisterBuffer_reg_4__6_ ( .D(queueRegister[46]), .CK(n551), 
        .Q(queueRegisterBuffer[46]) );
  DFFQX1TS queueRegisterBuffer_reg_4__7_ ( .D(queueRegister[47]), .CK(n551), 
        .Q(queueRegisterBuffer[47]) );
  DFFQX1TS queueRegisterBuffer_reg_4__8_ ( .D(queueRegister[48]), .CK(n552), 
        .Q(queueRegisterBuffer[48]) );
  DFFQX1TS queueRegisterBuffer_reg_0__9_ ( .D(queueRegister[9]), .CK(n544), 
        .Q(queueRegisterBuffer[9]) );
  DFFQX1TS queueRegisterBuffer_reg_0__0_ ( .D(queueRegister[0]), .CK(n545), 
        .Q(queueRegisterBuffer[0]) );
  DFFQX1TS queueRegisterBuffer_reg_0__1_ ( .D(queueRegister[1]), .CK(n545), 
        .Q(queueRegisterBuffer[1]) );
  DFFQX1TS queueRegisterBuffer_reg_0__2_ ( .D(queueRegister[2]), .CK(n545), 
        .Q(queueRegisterBuffer[2]) );
  DFFQX1TS queueRegisterBuffer_reg_0__3_ ( .D(queueRegister[3]), .CK(n545), 
        .Q(queueRegisterBuffer[3]) );
  DFFQX1TS queueRegisterBuffer_reg_0__4_ ( .D(queueRegister[4]), .CK(n546), 
        .Q(queueRegisterBuffer[4]) );
  DFFQX1TS queueRegisterBuffer_reg_0__5_ ( .D(queueRegister[5]), .CK(n546), 
        .Q(queueRegisterBuffer[5]) );
  DFFQX1TS queueRegisterBuffer_reg_0__6_ ( .D(queueRegister[6]), .CK(n546), 
        .Q(queueRegisterBuffer[6]) );
  DFFQX1TS queueRegisterBuffer_reg_0__7_ ( .D(queueRegister[7]), .CK(n546), 
        .Q(queueRegisterBuffer[7]) );
  DFFQX1TS queueRegisterBuffer_reg_0__8_ ( .D(queueRegister[8]), .CK(n547), 
        .Q(queueRegisterBuffer[8]) );
  DFFQX1TS queueRegisterBuffer_reg_1__9_ ( .D(queueRegister[19]), .CK(n539), 
        .Q(queueRegisterBuffer[19]) );
  DFFQX1TS queueRegisterBuffer_reg_1__0_ ( .D(queueRegister[10]), .CK(n540), 
        .Q(queueRegisterBuffer[10]) );
  DFFQX1TS queueRegisterBuffer_reg_1__1_ ( .D(queueRegister[11]), .CK(n540), 
        .Q(queueRegisterBuffer[11]) );
  DFFQX1TS queueRegisterBuffer_reg_1__2_ ( .D(queueRegister[12]), .CK(n540), 
        .Q(queueRegisterBuffer[12]) );
  DFFQX1TS queueRegisterBuffer_reg_1__3_ ( .D(queueRegister[13]), .CK(n540), 
        .Q(queueRegisterBuffer[13]) );
  DFFQX1TS queueRegisterBuffer_reg_1__4_ ( .D(queueRegister[14]), .CK(n541), 
        .Q(queueRegisterBuffer[14]) );
  DFFQX1TS queueRegisterBuffer_reg_1__5_ ( .D(queueRegister[15]), .CK(n541), 
        .Q(queueRegisterBuffer[15]) );
  DFFQX1TS queueRegisterBuffer_reg_1__6_ ( .D(queueRegister[16]), .CK(n541), 
        .Q(queueRegisterBuffer[16]) );
  DFFQX1TS queueRegisterBuffer_reg_1__7_ ( .D(queueRegister[17]), .CK(n541), 
        .Q(queueRegisterBuffer[17]) );
  DFFQX1TS queueRegisterBuffer_reg_1__8_ ( .D(queueRegister[18]), .CK(n542), 
        .Q(queueRegisterBuffer[18]) );
  DFFQX1TS queueRegisterBuffer_reg_2__9_ ( .D(queueRegister[29]), .CK(n547), 
        .Q(queueRegisterBuffer[29]) );
  DFFQX1TS queueRegisterBuffer_reg_2__0_ ( .D(queueRegister[20]), .CK(n547), 
        .Q(queueRegisterBuffer[20]) );
  DFFQX1TS queueRegisterBuffer_reg_2__1_ ( .D(queueRegister[21]), .CK(n547), 
        .Q(queueRegisterBuffer[21]) );
  DFFQX1TS queueRegisterBuffer_reg_2__2_ ( .D(queueRegister[22]), .CK(n548), 
        .Q(queueRegisterBuffer[22]) );
  DFFQX1TS queueRegisterBuffer_reg_2__3_ ( .D(queueRegister[23]), .CK(n548), 
        .Q(queueRegisterBuffer[23]) );
  DFFQX1TS queueRegisterBuffer_reg_2__4_ ( .D(queueRegister[24]), .CK(n548), 
        .Q(queueRegisterBuffer[24]) );
  DFFQX1TS queueRegisterBuffer_reg_2__5_ ( .D(queueRegister[25]), .CK(n548), 
        .Q(queueRegisterBuffer[25]) );
  DFFQX1TS queueRegisterBuffer_reg_2__6_ ( .D(queueRegister[26]), .CK(n549), 
        .Q(queueRegisterBuffer[26]) );
  DFFQX1TS queueRegisterBuffer_reg_2__7_ ( .D(queueRegister[27]), .CK(n549), 
        .Q(queueRegisterBuffer[27]) );
  DFFQX1TS queueRegisterBuffer_reg_2__8_ ( .D(queueRegister[28]), .CK(n549), 
        .Q(queueRegisterBuffer[28]) );
  DFFQX1TS queueRegisterBuffer_reg_3__9_ ( .D(queueRegister[39]), .CK(n537), 
        .Q(queueRegisterBuffer[39]) );
  DFFQX1TS queueRegisterBuffer_reg_3__0_ ( .D(queueRegister[30]), .CK(n537), 
        .Q(queueRegisterBuffer[30]) );
  DFFQX1TS queueRegisterBuffer_reg_3__1_ ( .D(queueRegister[31]), .CK(n537), 
        .Q(queueRegisterBuffer[31]) );
  DFFQX1TS queueRegisterBuffer_reg_3__2_ ( .D(queueRegister[32]), .CK(n538), 
        .Q(queueRegisterBuffer[32]) );
  DFFQX1TS queueRegisterBuffer_reg_3__3_ ( .D(queueRegister[33]), .CK(n538), 
        .Q(queueRegisterBuffer[33]) );
  DFFQX1TS queueRegisterBuffer_reg_3__4_ ( .D(queueRegister[34]), .CK(n538), 
        .Q(queueRegisterBuffer[34]) );
  DFFQX1TS queueRegisterBuffer_reg_3__5_ ( .D(queueRegister[35]), .CK(n538), 
        .Q(queueRegisterBuffer[35]) );
  DFFQX1TS queueRegisterBuffer_reg_3__6_ ( .D(queueRegister[36]), .CK(n539), 
        .Q(queueRegisterBuffer[36]) );
  DFFQX1TS queueRegisterBuffer_reg_3__7_ ( .D(queueRegister[37]), .CK(n539), 
        .Q(queueRegisterBuffer[37]) );
  DFFQX1TS queueRegisterBuffer_reg_3__8_ ( .D(queueRegister[38]), .CK(n539), 
        .Q(queueRegisterBuffer[38]) );
  DFFQX1TS queueRegisterBuffer_reg_6__3_ ( .D(queueRegister[63]), .CK(n519), 
        .Q(queueRegisterBuffer[63]) );
  DFFQX1TS queueRegisterBuffer_reg_6__6_ ( .D(queueRegister[66]), .CK(n515), 
        .Q(queueRegisterBuffer[66]) );
  DFFQX1TS queueRegisterBuffer_reg_6__8_ ( .D(queueRegister[68]), .CK(n515), 
        .Q(queueRegisterBuffer[68]) );
  DFFQX1TS queueRegisterBuffer_reg_6__2_ ( .D(queueRegister[62]), .CK(n517), 
        .Q(queueRegisterBuffer[62]) );
  DFFQX1TS queueRegisterBuffer_reg_6__4_ ( .D(queueRegister[64]), .CK(n516), 
        .Q(queueRegisterBuffer[64]) );
  DFFQX1TS queueRegisterBuffer_reg_6__5_ ( .D(queueRegister[65]), .CK(n520), 
        .Q(queueRegisterBuffer[65]) );
  DFFQX1TS queueRegisterBuffer_reg_6__7_ ( .D(queueRegister[67]), .CK(n518), 
        .Q(queueRegisterBuffer[67]) );
  DFFQX1TS queueRegisterBuffer_reg_6__9_ ( .D(queueRegister[69]), .CK(n552), 
        .Q(queueRegisterBuffer[69]) );
  DFFQX1TS queueRegisterBuffer_reg_6__0_ ( .D(queueRegister[60]), .CK(n552), 
        .Q(queueRegisterBuffer[60]) );
  DFFQX1TS queueRegisterBuffer_reg_6__1_ ( .D(queueRegister[61]), .CK(n552), 
        .Q(queueRegisterBuffer[61]) );
  DFFQX1TS queueEndPointerBuffer_reg_9_ ( .D(queueEndPointer[9]), .CK(n535), 
        .Q(queueEndPointerBuffer[9]) );
  DFFQX1TS queueEndPointerBuffer_reg_0_ ( .D(n246), .CK(n535), .Q(
        queueEndPointerBuffer[0]) );
  DFFQX1TS queueEndPointerBuffer_reg_4_ ( .D(queueEndPointer[4]), .CK(n536), 
        .Q(queueEndPointerBuffer[4]) );
  DFFQX1TS queueEndPointerBuffer_reg_7_ ( .D(queueEndPointer[7]), .CK(n537), 
        .Q(queueEndPointerBuffer[7]) );
  DFFQX1TS queueEndPointerBuffer_reg_1_ ( .D(queueEndPointer[1]), .CK(n535), 
        .Q(queueEndPointerBuffer[1]) );
  DFFQX1TS queueEndPointerBuffer_reg_2_ ( .D(n218), .CK(n535), .Q(
        queueEndPointerBuffer[2]) );
  DFFQX1TS queueEndPointerBuffer_reg_3_ ( .D(queueEndPointer[3]), .CK(n536), 
        .Q(queueEndPointerBuffer[3]) );
  DFFQX1TS queueEndPointerBuffer_reg_5_ ( .D(queueEndPointer[5]), .CK(n536), 
        .Q(queueEndPointerBuffer[5]) );
  DFFQX1TS queueEndPointerBuffer_reg_6_ ( .D(queueEndPointer[6]), .CK(n536), 
        .Q(queueEndPointerBuffer[6]) );
  DFFQX1TS queueEndPointerBuffer_reg_8_ ( .D(queueEndPointer[8]), .CK(n515), 
        .Q(queueEndPointerBuffer[8]) );
  TLATXLTS queueEmpty_reg ( .G(N126), .D(N127), .Q(queueEmpty) );
  DFFQX1TS queueRegister_reg_6__4_ ( .D(n133), .CK(clk), .Q(queueRegister[64])
         );
  DFFQX1TS queueRegister_reg_6__6_ ( .D(n119), .CK(clk), .Q(queueRegister[66])
         );
  DFFQX1TS queueRegister_reg_1__9_ ( .D(n173), .CK(clk), .Q(queueRegister[19])
         );
  DFFQX1TS queueRegister_reg_6__9_ ( .D(n168), .CK(clk), .Q(queueRegister[69])
         );
  DFFQX1TS queueRegister_reg_6__2_ ( .D(n147), .CK(clk), .Q(queueRegister[62])
         );
  DFFQX1TS queueRegister_reg_6__3_ ( .D(n140), .CK(clk), .Q(queueRegister[63])
         );
  DFFQX1TS queueRegister_reg_6__5_ ( .D(n1260), .CK(clk), .Q(queueRegister[65]) );
  DFFQX1TS queueRegister_reg_4__0_ ( .D(n163), .CK(clk), .Q(queueRegister[40])
         );
  DFFQX1TS queueRegister_reg_4__1_ ( .D(n156), .CK(clk), .Q(queueRegister[41])
         );
  DFFQX1TS queueRegister_reg_4__7_ ( .D(n114), .CK(clk), .Q(queueRegister[47])
         );
  DFFQX1TS queueRegister_reg_4__8_ ( .D(n1070), .CK(clk), .Q(queueRegister[48]) );
  DFFQX1TS queueRegister_reg_6__0_ ( .D(n161), .CK(clk), .Q(queueRegister[60])
         );
  DFFQX1TS queueRegister_reg_6__1_ ( .D(n154), .CK(clk), .Q(queueRegister[61])
         );
  DFFQX1TS queueRegister_reg_6__7_ ( .D(n112), .CK(clk), .Q(queueRegister[67])
         );
  DFFHQX8TS queueRegister_reg_3__9_ ( .D(n171), .CK(clk), .Q(queueRegister[39]) );
  DFFHQX8TS queueRegister_reg_2__9_ ( .D(n172), .CK(clk), .Q(queueRegister[29]) );
  DFFHQX8TS queueRegister_reg_3__4_ ( .D(n136), .CK(clk), .Q(queueRegister[34]) );
  DFFHQX8TS queueRegister_reg_2__3_ ( .D(n144), .CK(clk), .Q(queueRegister[23]) );
  DFFHQX8TS queueRegister_reg_2__4_ ( .D(n137), .CK(clk), .Q(queueRegister[24]) );
  DFFHQX8TS queueRegister_reg_2__6_ ( .D(n123), .CK(clk), .Q(queueRegister[26]) );
  DFFHQX8TS queueRegister_reg_3__3_ ( .D(n143), .CK(clk), .Q(queueRegister[33]) );
  DFFHQX8TS queueRegister_reg_2__5_ ( .D(n130), .CK(clk), .Q(queueRegister[25]) );
  DFFHQX8TS queueRegister_reg_3__1_ ( .D(n157), .CK(clk), .Q(queueRegister[31]) );
  DFFHQX8TS queueRegister_reg_3__7_ ( .D(n115), .CK(clk), .Q(queueRegister[37]) );
  DFFHQX8TS queueRegister_reg_2__0_ ( .D(n165), .CK(clk), .Q(queueRegister[20]) );
  DFFHQX8TS queueRegister_reg_2__1_ ( .D(n158), .CK(clk), .Q(queueRegister[21]) );
  DFFHQX8TS queueRegister_reg_2__7_ ( .D(n116), .CK(clk), .Q(queueRegister[27]) );
  DFFSX4TS queueEndPointer_reg_9_ ( .D(n512), .CK(clk), .SN(n484), .Q(n528), 
        .QN(queueEndPointer[9]) );
  DFFHQX8TS queueRegister_reg_2__8_ ( .D(n109), .CK(clk), .Q(queueRegister[28]) );
  DFFHQX8TS queueRegister_reg_2__2_ ( .D(n151), .CK(clk), .Q(queueRegister[22]) );
  DFFHQX8TS queueRegister_reg_3__2_ ( .D(n150), .CK(clk), .Q(queueRegister[32]) );
  DFFHQX8TS queueRegister_reg_5__4_ ( .D(n134), .CK(clk), .Q(queueRegister[54]) );
  DFFHQX8TS queueRegister_reg_5__6_ ( .D(n120), .CK(clk), .Q(queueRegister[56]) );
  DFFHQX8TS queueRegister_reg_0__2_ ( .D(n153), .CK(clk), .Q(queueRegister[2])
         );
  DFFHQX8TS queueRegister_reg_0__3_ ( .D(n146), .CK(clk), .Q(queueRegister[3])
         );
  DFFHQX8TS queueRegister_reg_0__4_ ( .D(n139), .CK(clk), .Q(queueRegister[4])
         );
  DFFHQX8TS queueRegister_reg_0__6_ ( .D(n125), .CK(clk), .Q(queueRegister[6])
         );
  DFFHQX8TS queueRegister_reg_5__3_ ( .D(n141), .CK(clk), .Q(queueRegister[53]) );
  DFFHQX8TS queueRegister_reg_0__9_ ( .D(n174), .CK(clk), .Q(queueRegister[9])
         );
  DFFHQX8TS queueRegister_reg_0__5_ ( .D(n132), .CK(clk), .Q(queueRegister[5])
         );
  DFFHQX8TS queueRegister_reg_4__9_ ( .D(n170), .CK(clk), .Q(queueRegister[49]) );
  DFFHQX8TS queueRegister_reg_5__0_ ( .D(n162), .CK(clk), .Q(queueRegister[50]) );
  DFFHQX8TS queueRegister_reg_5__1_ ( .D(n155), .CK(clk), .Q(queueRegister[51]) );
  DFFHQX8TS queueRegister_reg_5__8_ ( .D(n1060), .CK(clk), .Q(
        queueRegister[58]) );
  DFFHQX8TS queueRegister_reg_0__0_ ( .D(n167), .CK(clk), .Q(queueRegister[0])
         );
  DFFHQX8TS queueRegister_reg_0__1_ ( .D(n160), .CK(clk), .Q(queueRegister[1])
         );
  DFFHQX8TS queueRegister_reg_0__7_ ( .D(n118), .CK(clk), .Q(queueRegister[7])
         );
  DFFHQX8TS queueRegister_reg_0__8_ ( .D(n111), .CK(clk), .Q(queueRegister[8])
         );
  DFFNSRX1TS indexCounter_reg_9_ ( .D(n95), .CKN(clk), .SN(1'b1), .RN(n479), 
        .Q(indexCounter[9]), .QN(n514) );
  DFFHQX8TS queueRegister_reg_1__6_ ( .D(n124), .CK(clk), .Q(queueRegister[16]) );
  DFFHQX8TS queueRegister_reg_1__3_ ( .D(n145), .CK(clk), .Q(queueRegister[13]) );
  DFFHQX8TS queueRegister_reg_1__0_ ( .D(n166), .CK(clk), .Q(queueRegister[10]) );
  DFFHQX8TS queueRegister_reg_1__1_ ( .D(n159), .CK(clk), .Q(queueRegister[11]) );
  DFFHQX8TS queueRegister_reg_1__7_ ( .D(n117), .CK(clk), .Q(queueRegister[17]) );
  DFFHQX4TS queueRegister_reg_5__7_ ( .D(n113), .CK(clk), .Q(queueRegister[57]) );
  DFFHQX4TS queueRegister_reg_1__8_ ( .D(n110), .CK(clk), .Q(queueRegister[18]) );
  DFFHQX4TS queueRegister_reg_5__9_ ( .D(n169), .CK(clk), .Q(queueRegister[59]) );
  DFFHQX4TS queueRegister_reg_5__5_ ( .D(n1270), .CK(clk), .Q(
        queueRegister[55]) );
  DFFHQX4TS queueRegister_reg_4__5_ ( .D(n128), .CK(clk), .Q(queueRegister[45]) );
  DFFRHQX2TS queueEndPointer_reg_5_ ( .D(n178), .CK(clk), .RN(n219), .Q(
        queueEndPointer[5]) );
  DFFSHQX8TS queueEndPointer_reg_4_ ( .D(n513), .CK(clk), .SN(n220), .Q(n524)
         );
  DFFSX4TS queueEndPointer_reg_6_ ( .D(n475), .CK(clk), .SN(n220), .Q(n523), 
        .QN(queueEndPointer[6]) );
  DFFSX4TS queueEndPointer_reg_0_ ( .D(n215), .CK(clk), .SN(n219), .Q(n521), 
        .QN(queueEndPointer[0]) );
  DFFSHQX8TS queueEndPointer_reg_3_ ( .D(n498), .CK(clk), .SN(n219), .Q(n525)
         );
  DFFHQX8TS queueRegister_reg_3__8_ ( .D(n474), .CK(clk), .Q(queueRegister[38]) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_0_ ( .D(n94), .CKN(n477), .SN(1'b1), 
        .RN(n483), .Q(queueFrontPointerBuffer[0]), .QN(n508) );
  TLATXLTS finished_reg ( .G(N89), .D(N90), .Q(finished), .QN(n509) );
  DFFQX2TS queueRegister_reg_6__8_ ( .D(n1050), .CK(clk), .Q(queueRegister[68]) );
  DFFHQX4TS queueRegister_reg_3__6_ ( .D(n122), .CK(clk), .Q(queueRegister[36]) );
  DFFHQX4TS queueRegister_reg_3__5_ ( .D(n129), .CK(clk), .Q(queueRegister[35]) );
  DFFHQX4TS queueRegister_reg_3__0_ ( .D(n164), .CK(clk), .Q(queueRegister[30]) );
  DFFHQX4TS queueRegister_reg_4__4_ ( .D(n135), .CK(clk), .Q(queueRegister[44]) );
  DFFHQX4TS queueRegister_reg_4__6_ ( .D(n121), .CK(clk), .Q(queueRegister[46]) );
  DFFHQX4TS queueRegister_reg_5__2_ ( .D(n148), .CK(clk), .Q(queueRegister[52]) );
  DFFHQX4TS queueRegister_reg_4__2_ ( .D(n149), .CK(clk), .Q(queueRegister[42]) );
  DFFHQX4TS queueRegister_reg_4__3_ ( .D(n142), .CK(clk), .Q(queueRegister[43]) );
  DFFHQX4TS queueRegister_reg_1__4_ ( .D(n138), .CK(clk), .Q(queueRegister[14]) );
  DFFHQX4TS queueRegister_reg_1__2_ ( .D(n152), .CK(clk), .Q(queueRegister[12]) );
  DFFHQX4TS queueRegister_reg_1__5_ ( .D(n131), .CK(clk), .Q(queueRegister[15]) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_1_ ( .D(n93), .CKN(n485), .SN(1'b1), 
        .RN(n482), .Q(queueFrontPointerBuffer[1]), .QN(n496) );
  DFFRXLTS indexOut_reg_0_ ( .D(N107), .CK(n486), .RN(n489), .Q(indexOut[0])
         );
  DFFRXLTS indexOut_reg_1_ ( .D(N106), .CK(n485), .RN(n490), .Q(indexOut[1])
         );
  DFFRXLTS indexOut_reg_2_ ( .D(N105), .CK(n487), .RN(n491), .Q(indexOut[2])
         );
  DFFRXLTS indexOut_reg_3_ ( .D(N104), .CK(n488), .RN(n489), .Q(indexOut[3])
         );
  DFFRXLTS indexOut_reg_4_ ( .D(N103), .CK(n486), .RN(n490), .Q(indexOut[4])
         );
  DFFRXLTS indexOut_reg_5_ ( .D(N102), .CK(n485), .RN(n491), .Q(indexOut[5])
         );
  DFFRXLTS indexOut_reg_6_ ( .D(N101), .CK(n476), .RN(n489), .Q(indexOut[6])
         );
  DFFRXLTS indexOut_reg_7_ ( .D(N100), .CK(n488), .RN(n490), .Q(indexOut[7])
         );
  DFFRXLTS indexOut_reg_8_ ( .D(N99), .CK(n487), .RN(n491), .Q(indexOut[8]) );
  DFFRXLTS indexOut_reg_9_ ( .D(N98), .CK(n476), .RN(n489), .Q(indexOut[9]) );
  CLKMX2X2TS U201 ( .A(n446), .B(queueRegister[66]), .S0(n445), .Y(n119) );
  INVX4TS U202 ( .A(n212), .Y(n447) );
  NAND3X1TS U203 ( .A(n203), .B(n202), .C(n201), .Y(n200) );
  NAND2BXLTS U204 ( .AN(n372), .B(n185), .Y(n186) );
  OAI2BB1X2TS U205 ( .A0N(n199), .A1N(n259), .B0(n263), .Y(n195) );
  NOR3X1TS U206 ( .A(n261), .B(n262), .C(n259), .Y(n201) );
  NOR2BX1TS U207 ( .AN(n262), .B(n534), .Y(n249) );
  NAND2X4TS U208 ( .A(n214), .B(queueEndPointer[0]), .Y(n226) );
  AND2X2TS U209 ( .A(n261), .B(n238), .Y(n199) );
  NAND2BX1TS U210 ( .AN(n514), .B(n262), .Y(n263) );
  INVX4TS U211 ( .A(n405), .Y(n417) );
  INVX2TS U212 ( .A(n478), .Y(n408) );
  NAND2X2TS U213 ( .A(n525), .B(n524), .Y(n272) );
  OAI21XLTS U214 ( .A0(n256), .A1(n255), .B0(n254), .Y(n980) );
  MX2X2TS U215 ( .A(n458), .B(queueRegister[24]), .S0(n456), .Y(n137) );
  MX2X2TS U216 ( .A(n460), .B(queueRegister[64]), .S0(n459), .Y(n133) );
  XOR2X1TS U217 ( .A(n188), .B(n449), .Y(n256) );
  NAND2X2TS U218 ( .A(n193), .B(n260), .Y(n188) );
  CLKINVX6TS U219 ( .A(n521), .Y(n406) );
  NOR2X2TS U220 ( .A(n241), .B(n240), .Y(n270) );
  MX2X2TS U221 ( .A(n416), .B(queueRegister[65]), .S0(n277), .Y(n1260) );
  MX2X2TS U222 ( .A(n416), .B(queueRegister[5]), .S0(n421), .Y(n132) );
  MX2X2TS U223 ( .A(n416), .B(queueRegister[55]), .S0(n415), .Y(n1270) );
  MX2X2TS U224 ( .A(n444), .B(queueRegister[33]), .S0(n418), .Y(n143) );
  MX2X2TS U225 ( .A(n444), .B(queueRegister[23]), .S0(n456), .Y(n144) );
  MX2X2TS U226 ( .A(n444), .B(queueRegister[63]), .S0(n277), .Y(n140) );
  INVX6TS U227 ( .A(n405), .Y(n416) );
  NAND2X2TS U228 ( .A(n373), .B(n236), .Y(n278) );
  NAND2X6TS U229 ( .A(n443), .B(n442), .Y(n421) );
  NAND2X4TS U230 ( .A(n426), .B(n425), .Y(n415) );
  NOR2X8TS U231 ( .A(n245), .B(n211), .Y(n426) );
  XNOR2X1TS U232 ( .A(n193), .B(n458), .Y(n293) );
  CLKINVX6TS U233 ( .A(n277), .Y(n411) );
  BUFX12TS U234 ( .A(n424), .Y(n443) );
  CLKINVX3TS U235 ( .A(n529), .Y(n444) );
  CLKINVX3TS U236 ( .A(n530), .Y(n398) );
  MXI2X1TS U237 ( .A(n495), .B(n293), .S0(n509), .Y(n1000) );
  CLKINVX3TS U238 ( .A(n495), .Y(n458) );
  OAI21XLTS U239 ( .A0(n292), .A1(n185), .B0(n189), .Y(n990) );
  INVX6TS U240 ( .A(n433), .Y(n418) );
  CLKINVX6TS U241 ( .A(n226), .Y(n433) );
  CLKINVX3TS U242 ( .A(n453), .Y(n460) );
  CLKINVX2TS U243 ( .A(n509), .Y(n262) );
  INVX4TS U244 ( .A(n533), .Y(n192) );
  INVX2TS U245 ( .A(n509), .Y(n255) );
  NOR2X1TS U246 ( .A(n265), .B(n239), .Y(n221) );
  NOR2X1TS U247 ( .A(n478), .B(n526), .Y(n225) );
  NOR2X1TS U248 ( .A(n246), .B(n408), .Y(n423) );
  OR2X1TS U249 ( .A(queueEndPointer[4]), .B(n388), .Y(n266) );
  INVX2TS U250 ( .A(n238), .Y(n185) );
  CLKINVX3TS U251 ( .A(n410), .Y(n236) );
  INVX2TS U252 ( .A(n410), .Y(n432) );
  INVX2TS U253 ( .A(finished), .Y(n238) );
  OAI21XLTS U254 ( .A0(n187), .A1(n185), .B0(n186), .Y(n1010) );
  INVX4TS U255 ( .A(n411), .Y(n445) );
  CLKINVX2TS U256 ( .A(n531), .Y(n371) );
  INVX2TS U257 ( .A(n195), .Y(n198) );
  CLKINVX2TS U258 ( .A(n234), .Y(n235) );
  CLKINVX2TS U259 ( .A(n253), .Y(n254) );
  NOR2BX2TS U260 ( .AN(n185), .B(n532), .Y(n190) );
  INVX2TS U261 ( .A(n205), .Y(n202) );
  INVX2TS U262 ( .A(n204), .Y(n203) );
  NAND2BX2TS U263 ( .AN(n493), .B(n194), .Y(n204) );
  INVX2TS U264 ( .A(n278), .Y(n206) );
  CLKINVX1TS U265 ( .A(n239), .Y(n553) );
  INVX4TS U266 ( .A(n411), .Y(n459) );
  NAND4X1TS U267 ( .A(n200), .B(n197), .C(n198), .D(n196), .Y(n95) );
  INVX2TS U268 ( .A(n396), .Y(n437) );
  NAND2X2TS U269 ( .A(n199), .B(n204), .Y(n197) );
  NAND2X2TS U270 ( .A(n205), .B(n199), .Y(n196) );
  INVX2TS U271 ( .A(n190), .Y(n189) );
  NAND2X4TS U272 ( .A(n206), .B(n260), .Y(n205) );
  XNOR2X1TS U273 ( .A(n237), .B(n210), .Y(n187) );
  INVX4TS U274 ( .A(n211), .Y(n401) );
  CLKINVX2TS U275 ( .A(n391), .Y(n282) );
  INVX2TS U276 ( .A(n251), .Y(n449) );
  INVX3TS U277 ( .A(n251), .Y(n446) );
  INVX4TS U278 ( .A(n244), .Y(n405) );
  CLKINVX1TS U279 ( .A(n210), .Y(n372) );
  INVX2TS U280 ( .A(n525), .Y(queueEndPointer[3]) );
  INVX2TS U281 ( .A(n514), .Y(n261) );
  CLKBUFX2TS U282 ( .A(n461), .Y(n463) );
  OR2X2TS U283 ( .A(n523), .B(n393), .Y(n228) );
  OR2X2TS U284 ( .A(n394), .B(n393), .Y(n395) );
  INVX2TS U285 ( .A(n249), .Y(n250) );
  CLKINVX1TS U286 ( .A(n265), .Y(n388) );
  CLKBUFX2TS U287 ( .A(n328), .Y(n324) );
  INVX1TS U288 ( .A(n380), .Y(n381) );
  INVX1TS U289 ( .A(n439), .Y(n407) );
  INVX3TS U290 ( .A(n260), .Y(n207) );
  NAND2X1TS U291 ( .A(queueEndPointer[4]), .B(queueEndPointer[5]), .Y(n380) );
  INVX4TS U292 ( .A(n406), .Y(n288) );
  NOR2X4TS U293 ( .A(queueEndPointer[0]), .B(n218), .Y(n442) );
  INVX2TS U294 ( .A(n524), .Y(queueEndPointer[4]) );
  INVX1TS U295 ( .A(queueEndPointer[5]), .Y(n394) );
  INVX2TS U296 ( .A(n521), .Y(n246) );
  INVX2TS U297 ( .A(n499), .Y(n218) );
  INVX2TS U298 ( .A(indexCounter[0]), .Y(n412) );
  CLKINVX2TS U299 ( .A(n531), .Y(n419) );
  INVX1TS U300 ( .A(n239), .Y(n220) );
  INVX1TS U301 ( .A(n239), .Y(n219) );
  BUFX3TS U302 ( .A(resetInputQueue), .Y(n239) );
  CLKINVX6TS U303 ( .A(n289), .Y(n193) );
  NAND4X4TS U304 ( .A(n193), .B(n260), .C(n446), .D(n232), .Y(n233) );
  OAI21X2TS U305 ( .A0(n208), .A1(n262), .B0(n250), .Y(n97) );
  OAI21X2TS U306 ( .A0(n191), .A1(n255), .B0(n235), .Y(n96) );
  XOR2X4TS U307 ( .A(n233), .B(n192), .Y(n191) );
  XOR2X4TS U308 ( .A(n209), .B(n534), .Y(n208) );
  CLKBUFX2TS U309 ( .A(n257), .Y(n194) );
  AND2X8TS U310 ( .A(n244), .B(indexCounter[4]), .Y(n260) );
  NAND3X8TS U311 ( .A(n257), .B(n431), .C(n373), .Y(n289) );
  NOR3X4TS U312 ( .A(n207), .B(n289), .C(n493), .Y(n209) );
  INVX2TS U313 ( .A(n265), .Y(n393) );
  NAND2BX1TS U314 ( .AN(n437), .B(n528), .Y(n284) );
  NOR2X4TS U315 ( .A(n224), .B(n269), .Y(n276) );
  OR2X4TS U316 ( .A(n272), .B(n241), .Y(n224) );
  INVX2TS U317 ( .A(n287), .Y(n377) );
  MX2X1TS U318 ( .A(n409), .B(queueRegister[68]), .S0(n445), .Y(n1050) );
  XOR2XLTS U319 ( .A(n227), .B(n523), .Y(n229) );
  CLKMX2X2TS U320 ( .A(n417), .B(queueRegister[45]), .S0(n413), .Y(n128) );
  MX2X1TS U321 ( .A(n427), .B(queueRegister[18]), .S0(n402), .Y(n110) );
  MX2X1TS U322 ( .A(n399), .B(queueRegister[17]), .S0(n403), .Y(n117) );
  MX2X1TS U323 ( .A(n431), .B(queueRegister[11]), .S0(n454), .Y(n159) );
  MX2X1TS U324 ( .A(n417), .B(queueRegister[15]), .S0(n454), .Y(n131) );
  MX2X1TS U325 ( .A(n419), .B(queueRegister[12]), .S0(n403), .Y(n152) );
  MX2X1TS U326 ( .A(n460), .B(queueRegister[14]), .S0(n454), .Y(n138) );
  MX2X1TS U327 ( .A(n236), .B(queueRegister[51]), .S0(n448), .Y(n155) );
  MX2X1TS U328 ( .A(n414), .B(queueRegister[43]), .S0(n457), .Y(n142) );
  MX2X1TS U329 ( .A(n371), .B(queueRegister[42]), .S0(n413), .Y(n149) );
  MX2X1TS U330 ( .A(n419), .B(queueRegister[52]), .S0(n415), .Y(n148) );
  MX2X1TS U331 ( .A(n446), .B(queueRegister[46]), .S0(n457), .Y(n121) );
  MX2X1TS U332 ( .A(n458), .B(queueRegister[44]), .S0(n457), .Y(n135) );
  CLKMX2X2TS U333 ( .A(n460), .B(queueRegister[4]), .S0(n420), .Y(n139) );
  MX2X1TS U334 ( .A(n460), .B(queueRegister[54]), .S0(n455), .Y(n134) );
  MX2X1TS U335 ( .A(n435), .B(queueRegister[30]), .S0(n226), .Y(n164) );
  MX2X1TS U336 ( .A(n416), .B(queueRegister[35]), .S0(n418), .Y(n129) );
  MX2X1TS U337 ( .A(n449), .B(queueRegister[36]), .S0(n226), .Y(n122) );
  MX2X1TS U338 ( .A(n451), .B(queueRegister[62]), .S0(n459), .Y(n147) );
  MX2X1TS U339 ( .A(n286), .B(queueRegister[19]), .S0(n274), .Y(n173) );
  NAND2BX1TS U340 ( .AN(n437), .B(n522), .Y(n384) );
  OR2X1TS U341 ( .A(queueEndPointer[8]), .B(n388), .Y(n389) );
  XOR2X1TS U342 ( .A(n436), .B(queueEndPointer[0]), .Y(n438) );
  XOR2XLTS U343 ( .A(n398), .B(n238), .Y(n1040) );
  XOR2X1TS U344 ( .A(n371), .B(n278), .Y(n279) );
  NOR2BX1TS U345 ( .AN(finished), .B(n533), .Y(n234) );
  NOR2BX1TS U346 ( .AN(n255), .B(n251), .Y(n253) );
  NOR2X2TS U347 ( .A(n278), .B(n404), .Y(n237) );
  NOR2X8TS U348 ( .A(n245), .B(n211), .Y(n424) );
  INVX6TS U349 ( .A(n212), .Y(n429) );
  AND2X8TS U350 ( .A(n214), .B(n288), .Y(n212) );
  CLKBUFX2TS U351 ( .A(indexCounter[3]), .Y(n210) );
  BUFX8TS U352 ( .A(n269), .Y(n211) );
  CLKINVX1TS U353 ( .A(n251), .Y(n252) );
  INVX2TS U354 ( .A(n453), .Y(n290) );
  CLKINVX6TS U355 ( .A(n412), .Y(n373) );
  CLKBUFX2TS U356 ( .A(indexCounter[2]), .Y(n451) );
  INVX2TS U357 ( .A(n422), .Y(n399) );
  INVX2TS U358 ( .A(n437), .Y(n385) );
  INVX2TS U359 ( .A(n422), .Y(n434) );
  INVX2TS U360 ( .A(n422), .Y(n232) );
  XOR2X1TS U361 ( .A(n499), .B(n407), .Y(n213) );
  AND2X8TS U362 ( .A(n276), .B(n225), .Y(n214) );
  INVX4TS U363 ( .A(n433), .Y(n452) );
  XNOR2X1TS U364 ( .A(n246), .B(n393), .Y(n215) );
  OR2X1TS U365 ( .A(n500), .B(n496), .Y(n216) );
  OR2X1TS U366 ( .A(resetBuffer), .B(n515), .Y(n217) );
  NOR2XLTS U367 ( .A(queueFrontPointerBuffer[2]), .B(n496), .Y(n294) );
  NOR2XLTS U368 ( .A(n295), .B(n500), .Y(n296) );
  INVX2TS U369 ( .A(indexCounter[8]), .Y(n258) );
  INVX2TS U370 ( .A(n258), .Y(n427) );
  NAND2BX2TS U371 ( .AN(n255), .B(pixelValue), .Y(n265) );
  NAND2X2TS U372 ( .A(n523), .B(n221), .Y(n241) );
  NOR2X4TS U373 ( .A(queueEndPointer[9]), .B(queueEndPointer[8]), .Y(n223) );
  NOR2X4TS U374 ( .A(queueEndPointer[7]), .B(queueEndPointer[5]), .Y(n222) );
  NAND2X4TS U375 ( .A(n223), .B(n222), .Y(n269) );
  CLKMX2X2TS U376 ( .A(queueRegister[38]), .B(n427), .S0(n433), .Y(n474) );
  NAND4X2TS U377 ( .A(n406), .B(queueEndPointer[3]), .C(queueEndPointer[1]), 
        .D(n478), .Y(n391) );
  NOR2X1TS U378 ( .A(n391), .B(n380), .Y(n227) );
  INVX2TS U379 ( .A(n393), .Y(n396) );
  OAI21X1TS U380 ( .A0(n229), .A1(n396), .B0(n228), .Y(n230) );
  CLKINVX1TS U381 ( .A(n230), .Y(n475) );
  NAND2X2TS U382 ( .A(indexCounter[2]), .B(indexCounter[3]), .Y(n231) );
  CLKINVX6TS U383 ( .A(n231), .Y(n257) );
  INVX2TS U384 ( .A(indexCounter[1]), .Y(n410) );
  CLKINVX6TS U385 ( .A(n410), .Y(n431) );
  BUFX4TS U386 ( .A(indexCounter[5]), .Y(n244) );
  INVX2TS U387 ( .A(indexCounter[6]), .Y(n251) );
  INVX2TS U388 ( .A(indexCounter[7]), .Y(n422) );
  INVX2TS U389 ( .A(n258), .Y(n430) );
  INVX2TS U390 ( .A(n451), .Y(n404) );
  INVX2TS U391 ( .A(indexCounter[4]), .Y(n453) );
  INVX2TS U392 ( .A(n526), .Y(n240) );
  NAND2BX4TS U393 ( .AN(n272), .B(n270), .Y(n245) );
  NAND2X4TS U394 ( .A(n443), .B(n442), .Y(n420) );
  INVX2TS U395 ( .A(dequeue), .Y(n247) );
  INVX2TS U396 ( .A(n247), .Y(n487) );
  INVX2TS U397 ( .A(n487), .Y(n242) );
  INVX2TS U398 ( .A(n242), .Y(n476) );
  INVX2TS U399 ( .A(n242), .Y(n477) );
  INVX2TS U400 ( .A(n243), .Y(n484) );
  INVX2TS U401 ( .A(n553), .Y(n243) );
  INVX2TS U402 ( .A(n243), .Y(n479) );
  INVX2TS U403 ( .A(n243), .Y(n480) );
  NAND2X2TS U404 ( .A(n426), .B(n423), .Y(n413) );
  CLKBUFX2TS U405 ( .A(writeBufferEnable), .Y(n515) );
  INVX2TS U406 ( .A(n217), .Y(n481) );
  INVX2TS U407 ( .A(n217), .Y(n482) );
  INVX2TS U408 ( .A(n217), .Y(n483) );
  INVX2TS U409 ( .A(n247), .Y(n485) );
  INVX2TS U410 ( .A(n247), .Y(n486) );
  INVX2TS U411 ( .A(n247), .Y(n488) );
  CLKBUFX2TS U412 ( .A(resetBuffer), .Y(n248) );
  INVX2TS U413 ( .A(n248), .Y(n489) );
  INVX2TS U414 ( .A(n248), .Y(n490) );
  INVX2TS U415 ( .A(n248), .Y(n491) );
  INVX2TS U417 ( .A(n258), .Y(n409) );
  NAND2X2TS U418 ( .A(n399), .B(n409), .Y(n259) );
  CLKINVX1TS U419 ( .A(n282), .Y(n264) );
  XOR2X1TS U420 ( .A(n264), .B(n524), .Y(n267) );
  OAI21X1TS U421 ( .A0(n267), .A1(n265), .B0(n266), .Y(n513) );
  XNOR2X1TS U422 ( .A(n236), .B(n398), .Y(n268) );
  MXI2X1TS U423 ( .A(n268), .B(n494), .S0(finished), .Y(n1030) );
  INVX2TS U424 ( .A(indexCounter[9]), .Y(n287) );
  INVX2TS U425 ( .A(n287), .Y(n286) );
  NOR2X2TS U426 ( .A(n478), .B(n288), .Y(n271) );
  NAND2X2TS U427 ( .A(n271), .B(n270), .Y(n273) );
  NOR2X4TS U428 ( .A(n273), .B(n272), .Y(n400) );
  NAND2X1TS U429 ( .A(n401), .B(n400), .Y(n274) );
  NOR3X2TS U430 ( .A(n406), .B(n408), .C(n526), .Y(n275) );
  NAND2X4TS U431 ( .A(n276), .B(n275), .Y(n277) );
  CLKMX2X2TS U432 ( .A(n286), .B(queueRegister[69]), .S0(n445), .Y(n168) );
  MXI2X1TS U433 ( .A(n279), .B(n404), .S0(finished), .Y(n1020) );
  NAND2X1TS U434 ( .A(queueEndPointer[7]), .B(queueEndPointer[6]), .Y(n280) );
  NOR2X1TS U435 ( .A(n380), .B(n280), .Y(n281) );
  NAND2X2TS U436 ( .A(n282), .B(n281), .Y(n387) );
  NOR2X2TS U437 ( .A(n387), .B(n527), .Y(n283) );
  XNOR2X1TS U438 ( .A(n283), .B(n528), .Y(n285) );
  OAI21X1TS U439 ( .A0(n285), .A1(n385), .B0(n284), .Y(n512) );
  CLKMX2X2TS U440 ( .A(n286), .B(queueRegister[9]), .S0(n421), .Y(n174) );
  NOR2X2TS U441 ( .A(n288), .B(n408), .Y(n425) );
  CLKMX2X2TS U442 ( .A(n286), .B(queueRegister[59]), .S0(n415), .Y(n169) );
  CLKMX2X2TS U443 ( .A(n377), .B(queueRegister[49]), .S0(n413), .Y(n170) );
  CLKMX2X2TS U444 ( .A(n377), .B(queueRegister[29]), .S0(n429), .Y(n172) );
  CLKMX2X2TS U445 ( .A(n377), .B(queueRegister[39]), .S0(n418), .Y(n171) );
  NOR2BX2TS U446 ( .AN(n290), .B(n289), .Y(n291) );
  XOR2X1TS U447 ( .A(n291), .B(n532), .Y(n292) );
  INVX2TS U448 ( .A(n294), .Y(n304) );
  INVX2TS U449 ( .A(n304), .Y(n362) );
  OR2X1TS U450 ( .A(queueFrontPointerBuffer[2]), .B(queueFrontPointerBuffer[1]), .Y(n303) );
  INVX2TS U451 ( .A(n303), .Y(n363) );
  INVX2TS U452 ( .A(n496), .Y(n295) );
  INVX2TS U453 ( .A(n296), .Y(n305) );
  INVX2TS U454 ( .A(n305), .Y(n360) );
  AOI222XLTS U455 ( .A0(n362), .A1(queueRegisterBuffer[35]), .B0(n363), .B1(
        queueRegisterBuffer[15]), .C0(n360), .C1(queueRegisterBuffer[55]), .Y(
        n299) );
  INVX2TS U456 ( .A(n508), .Y(n310) );
  INVX2TS U457 ( .A(n310), .Y(n462) );
  INVX2TS U458 ( .A(n216), .Y(n335) );
  INVX2TS U459 ( .A(queueFrontPointerBuffer[0]), .Y(n311) );
  INVX2TS U460 ( .A(n311), .Y(n320) );
  INVX2TS U461 ( .A(n304), .Y(n330) );
  INVX2TS U462 ( .A(n303), .Y(n338) );
  INVX2TS U463 ( .A(n338), .Y(n309) );
  INVX2TS U464 ( .A(n309), .Y(n332) );
  INVX2TS U465 ( .A(n305), .Y(n328) );
  AOI222XLTS U466 ( .A0(n330), .A1(queueRegisterBuffer[25]), .B0(n332), .B1(
        queueRegisterBuffer[5]), .C0(n328), .C1(queueRegisterBuffer[45]), .Y(
        n297) );
  AOI2BB2XLTS U467 ( .B0(n335), .B1(queueRegisterBuffer[65]), .A0N(n320), 
        .A1N(n297), .Y(n298) );
  OAI21XLTS U468 ( .A0(n299), .A1(n462), .B0(n298), .Y(N102) );
  INVX2TS U469 ( .A(n304), .Y(n333) );
  INVX2TS U470 ( .A(n303), .Y(n340) );
  INVX2TS U471 ( .A(n305), .Y(n331) );
  AOI222XLTS U472 ( .A0(n333), .A1(queueRegisterBuffer[37]), .B0(n340), .B1(
        queueRegisterBuffer[17]), .C0(n331), .C1(queueRegisterBuffer[57]), .Y(
        n302) );
  INVX2TS U473 ( .A(n311), .Y(n366) );
  INVX2TS U474 ( .A(n330), .Y(n323) );
  INVX2TS U475 ( .A(n323), .Y(n318) );
  AOI222XLTS U476 ( .A0(n318), .A1(queueRegisterBuffer[27]), .B0(n340), .B1(
        queueRegisterBuffer[7]), .C0(n324), .C1(queueRegisterBuffer[47]), .Y(
        n300) );
  AOI2BB2XLTS U477 ( .B0(n335), .B1(queueRegisterBuffer[67]), .A0N(n366), 
        .A1N(n300), .Y(n301) );
  OAI21XLTS U478 ( .A0(n302), .A1(n462), .B0(n301), .Y(N100) );
  INVX2TS U479 ( .A(n303), .Y(n361) );
  AOI222XLTS U480 ( .A0(n330), .A1(queueRegisterBuffer[38]), .B0(n361), .B1(
        queueRegisterBuffer[18]), .C0(n328), .C1(queueRegisterBuffer[58]), .Y(
        n308) );
  INVX2TS U481 ( .A(n216), .Y(n367) );
  INVX2TS U482 ( .A(n305), .Y(n339) );
  AOI222XLTS U483 ( .A0(n294), .A1(queueRegisterBuffer[28]), .B0(n361), .B1(
        queueRegisterBuffer[8]), .C0(n339), .C1(queueRegisterBuffer[48]), .Y(
        n306) );
  AOI2BB2XLTS U484 ( .B0(n367), .B1(queueRegisterBuffer[68]), .A0N(n320), 
        .A1N(n306), .Y(n307) );
  OAI21XLTS U485 ( .A0(n308), .A1(n508), .B0(n307), .Y(N99) );
  INVX2TS U486 ( .A(n309), .Y(n329) );
  AOI222XLTS U487 ( .A0(n318), .A1(queueRegisterBuffer[33]), .B0(n329), .B1(
        queueRegisterBuffer[13]), .C0(n339), .C1(queueRegisterBuffer[53]), .Y(
        n314) );
  INVX2TS U488 ( .A(n310), .Y(n369) );
  AOI222XLTS U489 ( .A0(n362), .A1(queueRegisterBuffer[23]), .B0(n338), .B1(
        queueRegisterBuffer[3]), .C0(n360), .C1(queueRegisterBuffer[43]), .Y(
        n312) );
  AOI2BB2XLTS U490 ( .B0(n335), .B1(queueRegisterBuffer[63]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n312), .Y(n313) );
  OAI21XLTS U491 ( .A0(n314), .A1(n369), .B0(n313), .Y(N104) );
  AOI222XLTS U492 ( .A0(n362), .A1(queueRegisterBuffer[36]), .B0(n361), .B1(
        queueRegisterBuffer[16]), .C0(n360), .C1(queueRegisterBuffer[56]), .Y(
        n317) );
  AOI222XLTS U493 ( .A0(n333), .A1(queueRegisterBuffer[26]), .B0(n363), .B1(
        queueRegisterBuffer[6]), .C0(n331), .C1(queueRegisterBuffer[46]), .Y(
        n315) );
  AOI2BB2XLTS U494 ( .B0(n367), .B1(queueRegisterBuffer[66]), .A0N(n366), 
        .A1N(n315), .Y(n316) );
  OAI21XLTS U495 ( .A0(n317), .A1(n508), .B0(n316), .Y(N101) );
  AOI222XLTS U496 ( .A0(n318), .A1(queueRegisterBuffer[32]), .B0(n363), .B1(
        queueRegisterBuffer[12]), .C0(n324), .C1(queueRegisterBuffer[52]), .Y(
        n322) );
  AOI222XLTS U497 ( .A0(n333), .A1(queueRegisterBuffer[22]), .B0(n340), .B1(
        queueRegisterBuffer[2]), .C0(n331), .C1(queueRegisterBuffer[42]), .Y(
        n319) );
  AOI2BB2XLTS U498 ( .B0(n367), .B1(queueRegisterBuffer[62]), .A0N(n320), 
        .A1N(n319), .Y(n321) );
  OAI21XLTS U499 ( .A0(n322), .A1(n369), .B0(n321), .Y(N105) );
  AOI222XLTS U500 ( .A0(n294), .A1(queueRegisterBuffer[31]), .B0(n338), .B1(
        queueRegisterBuffer[11]), .C0(n339), .C1(queueRegisterBuffer[51]), .Y(
        n327) );
  INVX2TS U501 ( .A(n216), .Y(n465) );
  INVX2TS U502 ( .A(n323), .Y(n364) );
  AOI222XLTS U503 ( .A0(n364), .A1(queueRegisterBuffer[21]), .B0(n329), .B1(
        queueRegisterBuffer[1]), .C0(n324), .C1(queueRegisterBuffer[41]), .Y(
        n325) );
  AOI2BB2XLTS U504 ( .B0(n465), .B1(queueRegisterBuffer[61]), .A0N(n366), 
        .A1N(n325), .Y(n326) );
  OAI21XLTS U505 ( .A0(n327), .A1(n369), .B0(n326), .Y(N106) );
  AOI222XLTS U506 ( .A0(n330), .A1(queueRegisterBuffer[39]), .B0(n329), .B1(
        queueRegisterBuffer[19]), .C0(n328), .C1(queueRegisterBuffer[59]), .Y(
        n337) );
  AOI222XLTS U507 ( .A0(n333), .A1(queueRegisterBuffer[29]), .B0(n332), .B1(
        queueRegisterBuffer[9]), .C0(n331), .C1(queueRegisterBuffer[49]), .Y(
        n334) );
  AOI2BB2XLTS U508 ( .B0(n335), .B1(queueRegisterBuffer[69]), .A0N(n320), 
        .A1N(n334), .Y(n336) );
  OAI21XLTS U509 ( .A0(n337), .A1(n311), .B0(n336), .Y(N98) );
  AOI222XLTS U510 ( .A0(n364), .A1(queueRegisterBuffer[30]), .B0(n338), .B1(
        queueRegisterBuffer[10]), .C0(n296), .C1(queueRegisterBuffer[50]), .Y(
        n343) );
  AOI222XLTS U511 ( .A0(n318), .A1(queueRegisterBuffer[20]), .B0(n340), .B1(
        queueRegisterBuffer[0]), .C0(n339), .C1(queueRegisterBuffer[40]), .Y(
        n341) );
  AOI2BB2XLTS U512 ( .B0(n465), .B1(queueRegisterBuffer[60]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n341), .Y(n342) );
  OAI21XLTS U513 ( .A0(n343), .A1(n508), .B0(n342), .Y(N107) );
  XOR2XLTS U514 ( .A(n503), .B(queueEndPointerBuffer[3]), .Y(n345) );
  XOR2XLTS U515 ( .A(n500), .B(queueEndPointerBuffer[2]), .Y(n344) );
  NAND2X1TS U516 ( .A(n345), .B(n344), .Y(n359) );
  XOR2XLTS U517 ( .A(n502), .B(queueEndPointerBuffer[6]), .Y(n347) );
  XOR2XLTS U518 ( .A(n496), .B(queueEndPointerBuffer[1]), .Y(n346) );
  NAND2X1TS U519 ( .A(n347), .B(n346), .Y(n358) );
  XOR2XLTS U520 ( .A(n506), .B(queueEndPointerBuffer[8]), .Y(n349) );
  XOR2XLTS U521 ( .A(n507), .B(queueEndPointerBuffer[5]), .Y(n348) );
  NAND2X1TS U522 ( .A(n349), .B(n348), .Y(n357) );
  XNOR2X1TS U523 ( .A(n462), .B(queueEndPointerBuffer[0]), .Y(n351) );
  XNOR2X1TS U524 ( .A(n504), .B(queueEndPointerBuffer[9]), .Y(n350) );
  NOR2XLTS U525 ( .A(n351), .B(n350), .Y(n355) );
  XNOR2X1TS U526 ( .A(n501), .B(queueEndPointerBuffer[4]), .Y(n353) );
  XNOR2X1TS U527 ( .A(n505), .B(queueEndPointerBuffer[7]), .Y(n352) );
  NOR2XLTS U528 ( .A(n353), .B(n352), .Y(n354) );
  NAND3XLTS U529 ( .A(n481), .B(n355), .C(n354), .Y(n356) );
  NOR4XLTS U530 ( .A(n359), .B(n358), .C(n357), .D(n356), .Y(N127) );
  AOI222XLTS U531 ( .A0(n362), .A1(queueRegisterBuffer[34]), .B0(n361), .B1(
        queueRegisterBuffer[14]), .C0(n360), .C1(queueRegisterBuffer[54]), .Y(
        n370) );
  AOI222XLTS U532 ( .A0(n364), .A1(queueRegisterBuffer[24]), .B0(n363), .B1(
        queueRegisterBuffer[4]), .C0(n324), .C1(queueRegisterBuffer[44]), .Y(
        n365) );
  AOI2BB2XLTS U533 ( .B0(n367), .B1(queueRegisterBuffer[64]), .A0N(n366), 
        .A1N(n365), .Y(n368) );
  OAI21XLTS U534 ( .A0(n370), .A1(n369), .B0(n368), .Y(N103) );
  NAND4XLTS U535 ( .A(n371), .B(n534), .C(n493), .D(n484), .Y(n376) );
  NOR4XLTS U536 ( .A(n417), .B(n290), .C(n414), .D(n427), .Y(n374) );
  NAND3XLTS U537 ( .A(n431), .B(n374), .C(n530), .Y(n375) );
  NOR3XLTS U538 ( .A(n377), .B(n376), .C(n375), .Y(N90) );
  CLKBUFX2TS U539 ( .A(writeBufferEnable), .Y(n519) );
  CLKBUFX2TS U540 ( .A(n519), .Y(n520) );
  CLKBUFX2TS U541 ( .A(n520), .Y(n551) );
  CLKBUFX2TS U542 ( .A(n520), .Y(n550) );
  CLKBUFX2TS U543 ( .A(writeBufferEnable), .Y(n378) );
  CLKBUFX2TS U544 ( .A(n378), .Y(n544) );
  CLKBUFX2TS U545 ( .A(n378), .Y(n546) );
  CLKBUFX2TS U546 ( .A(n519), .Y(n379) );
  CLKBUFX2TS U547 ( .A(n379), .Y(n547) );
  CLKBUFX2TS U548 ( .A(n379), .Y(n548) );
  CLKBUFX2TS U549 ( .A(n379), .Y(n549) );
  CLKBUFX2TS U550 ( .A(n378), .Y(n545) );
  CLKBUFX2TS U551 ( .A(n378), .Y(n517) );
  CLKBUFX2TS U552 ( .A(n379), .Y(n518) );
  CLKBUFX2TS U553 ( .A(n520), .Y(n552) );
  CLKBUFX2TS U554 ( .A(n519), .Y(n516) );
  CLKBUFX2TS U555 ( .A(n516), .Y(n537) );
  CLKBUFX2TS U556 ( .A(n516), .Y(n535) );
  CLKBUFX2TS U557 ( .A(n516), .Y(n536) );
  NAND2X1TS U558 ( .A(n381), .B(queueEndPointer[6]), .Y(n382) );
  NOR2X1TS U559 ( .A(n382), .B(n391), .Y(n383) );
  XNOR2X1TS U560 ( .A(n383), .B(n522), .Y(n386) );
  OAI21X1TS U561 ( .A0(n386), .A1(n385), .B0(n384), .Y(n510) );
  XOR2X1TS U562 ( .A(n387), .B(n527), .Y(n390) );
  OAI21X1TS U563 ( .A0(n390), .A1(n385), .B0(n389), .Y(n511) );
  NOR2X1TS U564 ( .A(n391), .B(n524), .Y(n392) );
  XOR2X1TS U565 ( .A(n392), .B(n394), .Y(n397) );
  OAI21X1TS U566 ( .A0(n397), .A1(n396), .B0(n395), .Y(n178) );
  NAND2BXLTS U567 ( .AN(N90), .B(n480), .Y(N89) );
  CLKBUFX2TS U568 ( .A(n518), .Y(n543) );
  CLKBUFX2TS U569 ( .A(n517), .Y(n540) );
  CLKBUFX2TS U570 ( .A(n518), .Y(n541) );
  CLKBUFX2TS U571 ( .A(n518), .Y(n542) );
  CLKBUFX2TS U572 ( .A(n517), .Y(n538) );
  CLKBUFX2TS U573 ( .A(n517), .Y(n539) );
  NAND2X2TS U574 ( .A(n401), .B(n400), .Y(n403) );
  NAND2X2TS U575 ( .A(n401), .B(n400), .Y(n454) );
  CLKINVX1TS U576 ( .A(n529), .Y(n414) );
  CLKMX2X2TS U577 ( .A(n210), .B(queueRegister[13]), .S0(n403), .Y(n145) );
  NAND2X1TS U578 ( .A(n401), .B(n400), .Y(n402) );
  CLKINVX3TS U579 ( .A(n412), .Y(n435) );
  CLKMX2X2TS U580 ( .A(n435), .B(queueRegister[10]), .S0(n403), .Y(n166) );
  NAND2X1TS U581 ( .A(n406), .B(queueEndPointer[1]), .Y(n439) );
  MXI2X1TS U582 ( .A(n213), .B(n408), .S0(n396), .Y(n181) );
  CLKMX2X2TS U583 ( .A(n432), .B(queueRegister[61]), .S0(n459), .Y(n154) );
  CLKMX2X2TS U584 ( .A(n434), .B(queueRegister[67]), .S0(n445), .Y(n112) );
  CLKMX2X2TS U585 ( .A(n398), .B(queueRegister[60]), .S0(n459), .Y(n161) );
  NAND2X2TS U586 ( .A(n424), .B(n423), .Y(n457) );
  CLKMX2X2TS U587 ( .A(n210), .B(queueRegister[53]), .S0(n415), .Y(n141) );
  CLKMX2X2TS U588 ( .A(n417), .B(queueRegister[25]), .S0(n429), .Y(n130) );
  CLKMX2X2TS U589 ( .A(n419), .B(queueRegister[22]), .S0(n429), .Y(n151) );
  CLKMX2X2TS U590 ( .A(n419), .B(queueRegister[32]), .S0(n418), .Y(n150) );
  CLKMX2X2TS U591 ( .A(n430), .B(queueRegister[8]), .S0(n420), .Y(n111) );
  CLKMX2X2TS U592 ( .A(n434), .B(queueRegister[7]), .S0(n421), .Y(n118) );
  CLKMX2X2TS U593 ( .A(n432), .B(queueRegister[1]), .S0(n420), .Y(n160) );
  CLKMX2X2TS U594 ( .A(n373), .B(queueRegister[0]), .S0(n421), .Y(n167) );
  NAND2X2TS U595 ( .A(n426), .B(n425), .Y(n448) );
  CLKMX2X2TS U596 ( .A(n232), .B(queueRegister[57]), .S0(n448), .Y(n113) );
  NAND2X2TS U597 ( .A(n424), .B(n423), .Y(n428) );
  CLKMX2X2TS U598 ( .A(n432), .B(queueRegister[41]), .S0(n428), .Y(n156) );
  CLKMX2X2TS U599 ( .A(n430), .B(queueRegister[48]), .S0(n428), .Y(n1070) );
  NAND2X2TS U600 ( .A(n426), .B(n425), .Y(n455) );
  CLKMX2X2TS U601 ( .A(n427), .B(queueRegister[58]), .S0(n455), .Y(n1060) );
  CLKMX2X2TS U602 ( .A(n434), .B(queueRegister[47]), .S0(n428), .Y(n114) );
  CLKMX2X2TS U603 ( .A(n435), .B(queueRegister[40]), .S0(n457), .Y(n163) );
  CLKMX2X2TS U604 ( .A(n435), .B(queueRegister[50]), .S0(n455), .Y(n162) );
  CLKMX2X2TS U605 ( .A(n398), .B(queueRegister[20]), .S0(n429), .Y(n165) );
  CLKMX2X2TS U606 ( .A(n430), .B(queueRegister[28]), .S0(n447), .Y(n109) );
  INVX6TS U607 ( .A(n212), .Y(n456) );
  CLKMX2X2TS U608 ( .A(n431), .B(queueRegister[21]), .S0(n456), .Y(n158) );
  CLKMX2X2TS U609 ( .A(n232), .B(queueRegister[27]), .S0(n447), .Y(n116) );
  CLKMX2X2TS U610 ( .A(n236), .B(queueRegister[31]), .S0(n452), .Y(n157) );
  CLKMX2X2TS U611 ( .A(n434), .B(queueRegister[37]), .S0(n452), .Y(n115) );
  INVX2TS U612 ( .A(queueEndPointer[1]), .Y(n436) );
  CLKMX2X2TS U613 ( .A(n526), .B(n438), .S0(n437), .Y(n497) );
  NOR2X1TS U614 ( .A(n439), .B(n499), .Y(n440) );
  XNOR2X1TS U615 ( .A(n440), .B(n525), .Y(n441) );
  MXI2X1TS U616 ( .A(n441), .B(queueEndPointer[3]), .S0(n385), .Y(n498) );
  NAND2X4TS U617 ( .A(n443), .B(n442), .Y(n450) );
  CLKMX2X2TS U618 ( .A(n444), .B(queueRegister[3]), .S0(n450), .Y(n146) );
  CLKMX2X2TS U619 ( .A(n446), .B(queueRegister[6]), .S0(n450), .Y(n125) );
  CLKMX2X2TS U620 ( .A(n449), .B(queueRegister[26]), .S0(n447), .Y(n123) );
  CLKMX2X2TS U621 ( .A(n449), .B(queueRegister[56]), .S0(n448), .Y(n120) );
  CLKMX2X2TS U622 ( .A(n252), .B(queueRegister[16]), .S0(n454), .Y(n124) );
  CLKMX2X2TS U623 ( .A(n451), .B(queueRegister[2]), .S0(n450), .Y(n153) );
  CLKMX2X2TS U624 ( .A(n458), .B(queueRegister[34]), .S0(n452), .Y(n136) );
  NAND2BXLTS U625 ( .AN(N127), .B(n481), .Y(N126) );
  NOR2XLTS U626 ( .A(queueEmpty), .B(n311), .Y(n461) );
  AOI21X1TS U627 ( .A0(queueEmpty), .A1(n462), .B0(n461), .Y(n94) );
  AOI2BB2XLTS U628 ( .B0(queueFrontPointerBuffer[1]), .B1(n463), .A0N(n463), 
        .A1N(queueFrontPointerBuffer[1]), .Y(n93) );
  NAND2X1TS U629 ( .A(queueFrontPointerBuffer[1]), .B(n463), .Y(n464) );
  XNOR2X1TS U630 ( .A(queueFrontPointerBuffer[2]), .B(n464), .Y(n92) );
  NAND2X1TS U631 ( .A(n465), .B(n461), .Y(n467) );
  NAND3XLTS U632 ( .A(n465), .B(n463), .C(queueFrontPointerBuffer[3]), .Y(n468) );
  INVX2TS U633 ( .A(n468), .Y(n466) );
  AOI21X1TS U634 ( .A0(n467), .A1(n503), .B0(n466), .Y(n91) );
  NOR2XLTS U635 ( .A(n501), .B(n468), .Y(n469) );
  AOI21X1TS U636 ( .A0(n468), .A1(n501), .B0(n469), .Y(n900) );
  NAND2X1TS U637 ( .A(n469), .B(queueFrontPointerBuffer[5]), .Y(n470) );
  OA21XLTS U638 ( .A0(n469), .A1(queueFrontPointerBuffer[5]), .B0(n470), .Y(
        n890) );
  NOR2XLTS U639 ( .A(n502), .B(n470), .Y(n471) );
  AOI21X1TS U640 ( .A0(n470), .A1(n502), .B0(n471), .Y(n88) );
  NAND2X1TS U641 ( .A(n471), .B(queueFrontPointerBuffer[7]), .Y(n472) );
  OA21XLTS U642 ( .A0(n471), .A1(queueFrontPointerBuffer[7]), .B0(n472), .Y(
        n87) );
  XNOR2X1TS U643 ( .A(queueFrontPointerBuffer[8]), .B(n472), .Y(n86) );
  NAND2BXLTS U645 ( .AN(n472), .B(queueFrontPointerBuffer[8]), .Y(n473) );
  XNOR2X1TS U646 ( .A(queueFrontPointerBuffer[9]), .B(n473), .Y(n85) );
endmodule

