/*
 * This file describes the behaviour and IO of Layer 1. 
 * All modules needed for Layer 1 are instantiated here.
 */

`include "GlobalVariables.v"


module Layer1Controller (
	input clkIn,    // Clock
	input clk_en, // Clock Enable
	input reset,  // Asynchronous reset active low
	
);

endmodule