
module InputQueueRegister ( clk, resetInputQueue, resetBuffer, pixelValue, 
        dequeue, writeBufferEnable, finished, indexOut, queueEmpty );
  output [9:0] indexOut;
  input clk, resetInputQueue, resetBuffer, pixelValue, dequeue,
         writeBufferEnable;
  output finished, queueEmpty;
  wire   N89, N90, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N126, N127, n81, n83, n85, n86, n87, n88, n890, n900, n91, n92, n93,
         n94, n95, n96, n97, n980, n990, n1000, n1010, n1020, n1030, n1040,
         n1050, n1060, n1070, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n1260,
         n1270, n128, n129, n130, n131, n132, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n168, n169, n170, n171, n172,
         n173, n174, n181, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447;
  wire   [9:0] queueEndPointerBuffer;
  wire   [9:1] queueEndPointer;
  wire   [69:0] queueRegister;
  wire   [69:0] queueRegisterBuffer;
  wire   [9:0] indexCounter;
  wire   [9:0] queueFrontPointerBuffer;

  DFFNSRX1TS indexCounter_reg_6_ ( .D(n980), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[6]), .QN(n194) );
  DFFNSRX1TS indexCounter_reg_7_ ( .D(n97), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[7]), .QN(n445) );
  DFFNSRX1TS indexCounter_reg_8_ ( .D(n96), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[8]), .QN(n444) );
  DFFNSRX1TS indexCounter_reg_5_ ( .D(n990), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[5]), .QN(n443) );
  DFFNSRX1TS indexCounter_reg_2_ ( .D(n1020), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[2]), .QN(n441) );
  DFFNSRX1TS indexCounter_reg_3_ ( .D(n1010), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[3]), .QN(n439) );
  DFFNSRX1TS indexCounter_reg_9_ ( .D(n95), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[9]), .QN(n442) );
  DFFNSRX1TS indexCounter_reg_4_ ( .D(n1000), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[4]), .QN(n414) );
  DFFNSRX1TS indexCounter_reg_1_ ( .D(n1030), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[1]), .QN(n413) );
  DFFNSRX4TS indexCounter_reg_0_ ( .D(n1040), .CKN(clk), .SN(1'b1), .RN(n447), 
        .Q(indexCounter[0]), .QN(n440) );
  DFFSX4TS queueEndPointer_reg_1_ ( .D(n412), .CK(clk), .SN(n447), .Q(n436), 
        .QN(queueEndPointer[1]) );
  DFFSX4TS queueEndPointer_reg_7_ ( .D(n428), .CK(clk), .SN(n447), .Q(n431), 
        .QN(queueEndPointer[7]) );
  DFFSX4TS queueEndPointer_reg_3_ ( .D(n410), .CK(clk), .SN(n447), .Q(n434), 
        .QN(queueEndPointer[3]) );
  DFFSX4TS queueEndPointer_reg_9_ ( .D(n425), .CK(clk), .SN(n447), .Q(n438), 
        .QN(queueEndPointer[9]) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_0_ ( .D(n94), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[0]), .QN(n423) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_5_ ( .D(n890), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[5]), .QN(n422) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_8_ ( .D(n86), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[8]), .QN(n421) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_7_ ( .D(n87), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[7]), .QN(n420) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_9_ ( .D(n85), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[9]), .QN(n419) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_3_ ( .D(n91), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[3]), .QN(n418) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_6_ ( .D(n88), .CKN(n210), .SN(1'b1), 
        .RN(n83), .QN(n417) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_4_ ( .D(n900), .CKN(n210), .SN(1'b1), 
        .RN(n83), .QN(n416) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_2_ ( .D(n92), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[2]), .QN(n415) );
  DFFQX1TS queueRegisterBuffer_reg_5__9_ ( .D(queueRegister[59]), .CK(n429), 
        .Q(queueRegisterBuffer[59]) );
  DFFQX1TS queueRegisterBuffer_reg_5__0_ ( .D(queueRegister[50]), .CK(n429), 
        .Q(queueRegisterBuffer[50]) );
  DFFQX1TS queueRegisterBuffer_reg_5__1_ ( .D(queueRegister[51]), .CK(n429), 
        .Q(queueRegisterBuffer[51]) );
  DFFQX1TS queueRegisterBuffer_reg_5__2_ ( .D(queueRegister[52]), .CK(n429), 
        .Q(queueRegisterBuffer[52]) );
  DFFQX1TS queueRegisterBuffer_reg_5__3_ ( .D(queueRegister[53]), .CK(n429), 
        .Q(queueRegisterBuffer[53]) );
  DFFQX1TS queueRegisterBuffer_reg_5__4_ ( .D(queueRegister[54]), .CK(n429), 
        .Q(queueRegisterBuffer[54]) );
  DFFQX1TS queueRegisterBuffer_reg_5__5_ ( .D(queueRegister[55]), .CK(n429), 
        .Q(queueRegisterBuffer[55]) );
  DFFQX1TS queueRegisterBuffer_reg_5__6_ ( .D(queueRegister[56]), .CK(n429), 
        .Q(queueRegisterBuffer[56]) );
  DFFQX1TS queueRegisterBuffer_reg_5__7_ ( .D(queueRegister[57]), .CK(n429), 
        .Q(queueRegisterBuffer[57]) );
  DFFQX1TS queueRegisterBuffer_reg_5__8_ ( .D(queueRegister[58]), .CK(n429), 
        .Q(queueRegisterBuffer[58]) );
  DFFQX1TS queueRegisterBuffer_reg_4__9_ ( .D(queueRegister[49]), .CK(n429), 
        .Q(queueRegisterBuffer[49]) );
  DFFQX1TS queueRegisterBuffer_reg_4__0_ ( .D(queueRegister[40]), .CK(n429), 
        .Q(queueRegisterBuffer[40]) );
  DFFQX1TS queueRegisterBuffer_reg_4__1_ ( .D(queueRegister[41]), .CK(n429), 
        .Q(queueRegisterBuffer[41]) );
  DFFQX1TS queueRegisterBuffer_reg_4__2_ ( .D(queueRegister[42]), .CK(n429), 
        .Q(queueRegisterBuffer[42]) );
  DFFQX1TS queueRegisterBuffer_reg_4__3_ ( .D(queueRegister[43]), .CK(n429), 
        .Q(queueRegisterBuffer[43]) );
  DFFQX1TS queueRegisterBuffer_reg_4__4_ ( .D(queueRegister[44]), .CK(n429), 
        .Q(queueRegisterBuffer[44]) );
  DFFQX1TS queueRegisterBuffer_reg_4__5_ ( .D(queueRegister[45]), .CK(n429), 
        .Q(queueRegisterBuffer[45]) );
  DFFQX1TS queueRegisterBuffer_reg_4__6_ ( .D(queueRegister[46]), .CK(n429), 
        .Q(queueRegisterBuffer[46]) );
  DFFQX1TS queueRegisterBuffer_reg_4__7_ ( .D(queueRegister[47]), .CK(n429), 
        .Q(queueRegisterBuffer[47]) );
  DFFQX1TS queueRegisterBuffer_reg_4__8_ ( .D(queueRegister[48]), .CK(n429), 
        .Q(queueRegisterBuffer[48]) );
  DFFQX1TS queueRegisterBuffer_reg_1__9_ ( .D(queueRegister[19]), .CK(n429), 
        .Q(queueRegisterBuffer[19]) );
  DFFQX1TS queueRegisterBuffer_reg_1__0_ ( .D(queueRegister[10]), .CK(n429), 
        .Q(queueRegisterBuffer[10]) );
  DFFQX1TS queueRegisterBuffer_reg_1__1_ ( .D(queueRegister[11]), .CK(n429), 
        .Q(queueRegisterBuffer[11]) );
  DFFQX1TS queueRegisterBuffer_reg_1__2_ ( .D(queueRegister[12]), .CK(n429), 
        .Q(queueRegisterBuffer[12]) );
  DFFQX1TS queueRegisterBuffer_reg_1__3_ ( .D(queueRegister[13]), .CK(n429), 
        .Q(queueRegisterBuffer[13]) );
  DFFQX1TS queueRegisterBuffer_reg_1__4_ ( .D(queueRegister[14]), .CK(n429), 
        .Q(queueRegisterBuffer[14]) );
  DFFQX1TS queueRegisterBuffer_reg_1__5_ ( .D(queueRegister[15]), .CK(n429), 
        .Q(queueRegisterBuffer[15]) );
  DFFQX1TS queueRegisterBuffer_reg_1__6_ ( .D(queueRegister[16]), .CK(n429), 
        .Q(queueRegisterBuffer[16]) );
  DFFQX1TS queueRegisterBuffer_reg_1__7_ ( .D(queueRegister[17]), .CK(n429), 
        .Q(queueRegisterBuffer[17]) );
  DFFQX1TS queueRegisterBuffer_reg_1__8_ ( .D(queueRegister[18]), .CK(n429), 
        .Q(queueRegisterBuffer[18]) );
  DFFQX1TS queueRegisterBuffer_reg_0__9_ ( .D(queueRegister[9]), .CK(n429), 
        .Q(queueRegisterBuffer[9]) );
  DFFQX1TS queueRegisterBuffer_reg_0__0_ ( .D(queueRegister[0]), .CK(n429), 
        .Q(queueRegisterBuffer[0]) );
  DFFQX1TS queueRegisterBuffer_reg_0__1_ ( .D(queueRegister[1]), .CK(n429), 
        .Q(queueRegisterBuffer[1]) );
  DFFQX1TS queueRegisterBuffer_reg_0__2_ ( .D(queueRegister[2]), .CK(n429), 
        .Q(queueRegisterBuffer[2]) );
  DFFQX1TS queueRegisterBuffer_reg_0__3_ ( .D(queueRegister[3]), .CK(n429), 
        .Q(queueRegisterBuffer[3]) );
  DFFQX1TS queueRegisterBuffer_reg_0__4_ ( .D(queueRegister[4]), .CK(n429), 
        .Q(queueRegisterBuffer[4]) );
  DFFQX1TS queueRegisterBuffer_reg_0__5_ ( .D(queueRegister[5]), .CK(n429), 
        .Q(queueRegisterBuffer[5]) );
  DFFQX1TS queueRegisterBuffer_reg_0__6_ ( .D(queueRegister[6]), .CK(n429), 
        .Q(queueRegisterBuffer[6]) );
  DFFQX1TS queueRegisterBuffer_reg_0__7_ ( .D(queueRegister[7]), .CK(n429), 
        .Q(queueRegisterBuffer[7]) );
  DFFQX1TS queueRegisterBuffer_reg_0__8_ ( .D(queueRegister[8]), .CK(n429), 
        .Q(queueRegisterBuffer[8]) );
  DFFQX1TS queueRegisterBuffer_reg_3__9_ ( .D(queueRegister[39]), .CK(n429), 
        .Q(queueRegisterBuffer[39]) );
  DFFQX1TS queueRegisterBuffer_reg_3__0_ ( .D(queueRegister[30]), .CK(n429), 
        .Q(queueRegisterBuffer[30]) );
  DFFQX1TS queueRegisterBuffer_reg_3__1_ ( .D(queueRegister[31]), .CK(n429), 
        .Q(queueRegisterBuffer[31]) );
  DFFQX1TS queueRegisterBuffer_reg_3__2_ ( .D(queueRegister[32]), .CK(n429), 
        .Q(queueRegisterBuffer[32]) );
  DFFQX1TS queueRegisterBuffer_reg_3__3_ ( .D(queueRegister[33]), .CK(n429), 
        .Q(queueRegisterBuffer[33]) );
  DFFQX1TS queueRegisterBuffer_reg_3__4_ ( .D(queueRegister[34]), .CK(n429), 
        .Q(queueRegisterBuffer[34]) );
  DFFQX1TS queueRegisterBuffer_reg_3__5_ ( .D(queueRegister[35]), .CK(n429), 
        .Q(queueRegisterBuffer[35]) );
  DFFQX1TS queueRegisterBuffer_reg_3__6_ ( .D(queueRegister[36]), .CK(n429), 
        .Q(queueRegisterBuffer[36]) );
  DFFQX1TS queueRegisterBuffer_reg_3__7_ ( .D(queueRegister[37]), .CK(n429), 
        .Q(queueRegisterBuffer[37]) );
  DFFQX1TS queueRegisterBuffer_reg_3__8_ ( .D(queueRegister[38]), .CK(n429), 
        .Q(queueRegisterBuffer[38]) );
  DFFQX1TS queueRegisterBuffer_reg_2__9_ ( .D(queueRegister[29]), .CK(n429), 
        .Q(queueRegisterBuffer[29]) );
  DFFQX1TS queueRegisterBuffer_reg_2__0_ ( .D(queueRegister[20]), .CK(n429), 
        .Q(queueRegisterBuffer[20]) );
  DFFQX1TS queueRegisterBuffer_reg_2__1_ ( .D(queueRegister[21]), .CK(n429), 
        .Q(queueRegisterBuffer[21]) );
  DFFQX1TS queueRegisterBuffer_reg_2__2_ ( .D(queueRegister[22]), .CK(n429), 
        .Q(queueRegisterBuffer[22]) );
  DFFQX1TS queueRegisterBuffer_reg_2__3_ ( .D(queueRegister[23]), .CK(n429), 
        .Q(queueRegisterBuffer[23]) );
  DFFQX1TS queueRegisterBuffer_reg_2__4_ ( .D(queueRegister[24]), .CK(n429), 
        .Q(queueRegisterBuffer[24]) );
  DFFQX1TS queueRegisterBuffer_reg_2__5_ ( .D(queueRegister[25]), .CK(n429), 
        .Q(queueRegisterBuffer[25]) );
  DFFQX1TS queueRegisterBuffer_reg_2__6_ ( .D(queueRegister[26]), .CK(n429), 
        .Q(queueRegisterBuffer[26]) );
  DFFQX1TS queueRegisterBuffer_reg_2__7_ ( .D(queueRegister[27]), .CK(n429), 
        .Q(queueRegisterBuffer[27]) );
  DFFQX1TS queueRegisterBuffer_reg_2__8_ ( .D(queueRegister[28]), .CK(n429), 
        .Q(queueRegisterBuffer[28]) );
  DFFQX1TS queueRegisterBuffer_reg_6__9_ ( .D(queueRegister[69]), .CK(n429), 
        .Q(queueRegisterBuffer[69]) );
  DFFQX1TS queueRegisterBuffer_reg_6__0_ ( .D(queueRegister[60]), .CK(n429), 
        .Q(queueRegisterBuffer[60]) );
  DFFQX1TS queueRegisterBuffer_reg_6__1_ ( .D(queueRegister[61]), .CK(n429), 
        .Q(queueRegisterBuffer[61]) );
  DFFQX1TS queueRegisterBuffer_reg_6__2_ ( .D(queueRegister[62]), .CK(n429), 
        .Q(queueRegisterBuffer[62]) );
  DFFQX1TS queueRegisterBuffer_reg_6__3_ ( .D(queueRegister[63]), .CK(n429), 
        .Q(queueRegisterBuffer[63]) );
  DFFQX1TS queueRegisterBuffer_reg_6__4_ ( .D(queueRegister[64]), .CK(n429), 
        .Q(queueRegisterBuffer[64]) );
  DFFQX1TS queueRegisterBuffer_reg_6__5_ ( .D(queueRegister[65]), .CK(n429), 
        .Q(queueRegisterBuffer[65]) );
  DFFQX1TS queueRegisterBuffer_reg_6__6_ ( .D(queueRegister[66]), .CK(n429), 
        .Q(queueRegisterBuffer[66]) );
  DFFQX1TS queueRegisterBuffer_reg_6__7_ ( .D(queueRegister[67]), .CK(n429), 
        .Q(queueRegisterBuffer[67]) );
  DFFQX1TS queueRegisterBuffer_reg_6__8_ ( .D(queueRegister[68]), .CK(n429), 
        .Q(queueRegisterBuffer[68]) );
  DFFQX1TS queueEndPointerBuffer_reg_9_ ( .D(queueEndPointer[9]), .CK(n429), 
        .Q(queueEndPointerBuffer[9]) );
  DFFQX1TS queueEndPointerBuffer_reg_0_ ( .D(n446), .CK(n429), .Q(
        queueEndPointerBuffer[0]) );
  DFFQX1TS queueEndPointerBuffer_reg_4_ ( .D(queueEndPointer[4]), .CK(n429), 
        .Q(queueEndPointerBuffer[4]) );
  DFFQX1TS queueEndPointerBuffer_reg_1_ ( .D(queueEndPointer[1]), .CK(n429), 
        .Q(queueEndPointerBuffer[1]) );
  DFFQX1TS queueEndPointerBuffer_reg_2_ ( .D(queueEndPointer[2]), .CK(n429), 
        .Q(queueEndPointerBuffer[2]) );
  DFFQX1TS queueEndPointerBuffer_reg_3_ ( .D(queueEndPointer[3]), .CK(n429), 
        .Q(queueEndPointerBuffer[3]) );
  DFFQX1TS queueEndPointerBuffer_reg_5_ ( .D(queueEndPointer[5]), .CK(n429), 
        .Q(queueEndPointerBuffer[5]) );
  DFFQX1TS queueEndPointerBuffer_reg_6_ ( .D(queueEndPointer[6]), .CK(n429), 
        .Q(queueEndPointerBuffer[6]) );
  DFFQX1TS queueEndPointerBuffer_reg_8_ ( .D(queueEndPointer[8]), .CK(n429), 
        .Q(queueEndPointerBuffer[8]) );
  TLATXLTS queueEmpty_reg ( .G(N126), .D(N127), .Q(queueEmpty) );
  DFFRXLTS indexOut_reg_9_ ( .D(N98), .CK(n210), .RN(n81), .Q(indexOut[9]) );
  DFFRXLTS indexOut_reg_8_ ( .D(N99), .CK(n210), .RN(n81), .Q(indexOut[8]) );
  DFFRXLTS indexOut_reg_7_ ( .D(N100), .CK(n210), .RN(n81), .Q(indexOut[7]) );
  DFFRXLTS indexOut_reg_6_ ( .D(N101), .CK(n210), .RN(n81), .Q(indexOut[6]) );
  DFFRXLTS indexOut_reg_5_ ( .D(N102), .CK(n210), .RN(n81), .Q(indexOut[5]) );
  DFFRXLTS indexOut_reg_4_ ( .D(N103), .CK(n210), .RN(n81), .Q(indexOut[4]) );
  DFFRXLTS indexOut_reg_3_ ( .D(N104), .CK(n210), .RN(n81), .Q(indexOut[3]) );
  DFFRXLTS indexOut_reg_2_ ( .D(N105), .CK(n210), .RN(n81), .Q(indexOut[2]) );
  DFFRXLTS indexOut_reg_1_ ( .D(N106), .CK(n210), .RN(n81), .Q(indexOut[1]) );
  DFFRXLTS indexOut_reg_0_ ( .D(N107), .CK(n210), .RN(n81), .Q(indexOut[0]) );
  DFFQX1TS queueEndPointerBuffer_reg_7_ ( .D(queueEndPointer[7]), .CK(n429), 
        .Q(queueEndPointerBuffer[7]) );
  DFFQX1TS queueRegister_reg_0__4_ ( .D(n139), .CK(clk), .Q(queueRegister[4])
         );
  DFFQX1TS queueRegister_reg_0__6_ ( .D(n125), .CK(clk), .Q(queueRegister[6])
         );
  DFFQX1TS queueRegister_reg_2__4_ ( .D(n137), .CK(clk), .Q(queueRegister[24])
         );
  DFFQX1TS queueRegister_reg_2__6_ ( .D(n123), .CK(clk), .Q(queueRegister[26])
         );
  DFFQX1TS queueRegister_reg_0__9_ ( .D(n174), .CK(clk), .Q(queueRegister[9])
         );
  DFFQX1TS queueRegister_reg_0__2_ ( .D(n153), .CK(clk), .Q(queueRegister[2])
         );
  DFFQX1TS queueRegister_reg_0__5_ ( .D(n132), .CK(clk), .Q(queueRegister[5])
         );
  DFFQX1TS queueRegister_reg_2__9_ ( .D(n172), .CK(clk), .Q(queueRegister[29])
         );
  DFFQX1TS queueRegister_reg_2__5_ ( .D(n130), .CK(clk), .Q(queueRegister[25])
         );
  DFFQX1TS queueRegister_reg_3__0_ ( .D(n164), .CK(clk), .Q(queueRegister[30])
         );
  DFFQX1TS queueRegister_reg_0__1_ ( .D(n160), .CK(clk), .Q(queueRegister[1])
         );
  DFFQX1TS queueRegister_reg_0__7_ ( .D(n118), .CK(clk), .Q(queueRegister[7])
         );
  DFFQX1TS queueRegister_reg_2__7_ ( .D(n116), .CK(clk), .Q(queueRegister[27])
         );
  DFFQX1TS queueRegister_reg_2__8_ ( .D(n109), .CK(clk), .Q(queueRegister[28])
         );
  DFFHQX8TS queueRegister_reg_3__6_ ( .D(n122), .CK(clk), .Q(queueRegister[36]) );
  DFFHQX8TS queueRegister_reg_3__3_ ( .D(n143), .CK(clk), .Q(queueRegister[33]) );
  DFFHQX8TS queueRegister_reg_3__5_ ( .D(n129), .CK(clk), .Q(queueRegister[35]) );
  DFFHQX8TS queueRegister_reg_3__7_ ( .D(n115), .CK(clk), .Q(queueRegister[37]) );
  DFFHQX8TS queueRegister_reg_3__8_ ( .D(n108), .CK(clk), .Q(queueRegister[38]) );
  DFFHQX8TS queueRegister_reg_3__1_ ( .D(n157), .CK(clk), .Q(queueRegister[31]) );
  DFFHQX8TS queueRegister_reg_6__6_ ( .D(n119), .CK(clk), .Q(queueRegister[66]) );
  DFFHQX8TS queueRegister_reg_6__3_ ( .D(n140), .CK(clk), .Q(queueRegister[63]) );
  DFFHQX8TS queueRegister_reg_5__4_ ( .D(n134), .CK(clk), .Q(queueRegister[54]) );
  DFFHQX8TS queueRegister_reg_5__6_ ( .D(n120), .CK(clk), .Q(queueRegister[56]) );
  DFFHQX8TS queueRegister_reg_5__3_ ( .D(n141), .CK(clk), .Q(queueRegister[53]) );
  DFFHQX8TS queueRegister_reg_5__5_ ( .D(n1270), .CK(clk), .Q(
        queueRegister[55]) );
  DFFHQX8TS queueRegister_reg_5__1_ ( .D(n155), .CK(clk), .Q(queueRegister[51]) );
  DFFHQX8TS queueRegister_reg_5__7_ ( .D(n113), .CK(clk), .Q(queueRegister[57]) );
  DFFHQX8TS queueRegister_reg_5__8_ ( .D(n1060), .CK(clk), .Q(
        queueRegister[58]) );
  DFFHQX4TS queueRegister_reg_0__3_ ( .D(n146), .CK(clk), .Q(queueRegister[3])
         );
  DFFHQX4TS queueRegister_reg_2__3_ ( .D(n144), .CK(clk), .Q(queueRegister[23]) );
  DFFHQX4TS queueRegister_reg_1__3_ ( .D(n145), .CK(clk), .Q(queueRegister[13]) );
  DFFHQX4TS queueRegister_reg_4__3_ ( .D(n142), .CK(clk), .Q(queueRegister[43]) );
  DFFHQX4TS queueRegister_reg_1__2_ ( .D(n152), .CK(clk), .Q(queueRegister[12]) );
  DFFHQX4TS queueRegister_reg_2__2_ ( .D(n151), .CK(clk), .Q(queueRegister[22]) );
  DFFX4TS queueRegister_reg_5__0_ ( .D(n162), .CK(clk), .Q(queueRegister[50])
         );
  DFFX4TS queueRegister_reg_6__0_ ( .D(n161), .CK(clk), .Q(queueRegister[60])
         );
  DFFX4TS queueRegister_reg_2__0_ ( .D(n165), .CK(clk), .Q(queueRegister[20])
         );
  DFFHQX8TS queueRegister_reg_4__1_ ( .D(n156), .CK(clk), .Q(queueRegister[41]) );
  DFFHQX8TS queueRegister_reg_1__5_ ( .D(n131), .CK(clk), .Q(queueRegister[15]) );
  DFFHQX4TS queueRegister_reg_1__9_ ( .D(n173), .CK(clk), .Q(queueRegister[19]) );
  DFFHQX8TS queueRegister_reg_4__6_ ( .D(n121), .CK(clk), .Q(queueRegister[46]) );
  DFFHQX8TS queueRegister_reg_4__4_ ( .D(n135), .CK(clk), .Q(queueRegister[44]) );
  DFFHQX8TS queueRegister_reg_1__6_ ( .D(n124), .CK(clk), .Q(queueRegister[16]) );
  DFFHQX8TS queueRegister_reg_1__4_ ( .D(n138), .CK(clk), .Q(queueRegister[14]) );
  DFFHQX8TS queueRegister_reg_4__8_ ( .D(n1070), .CK(clk), .Q(
        queueRegister[48]) );
  DFFHQX8TS queueRegister_reg_4__7_ ( .D(n114), .CK(clk), .Q(queueRegister[47]) );
  DFFHQX8TS queueRegister_reg_4__2_ ( .D(n149), .CK(clk), .Q(queueRegister[42]) );
  DFFHQX4TS queueRegister_reg_4__9_ ( .D(n170), .CK(clk), .Q(queueRegister[49]) );
  DFFHQX8TS queueRegister_reg_1__1_ ( .D(n159), .CK(clk), .Q(queueRegister[11]) );
  DFFHQX8TS queueRegister_reg_4__5_ ( .D(n128), .CK(clk), .Q(queueRegister[45]) );
  DFFHQX8TS queueRegister_reg_1__7_ ( .D(n117), .CK(clk), .Q(queueRegister[17]) );
  DFFHQX8TS queueRegister_reg_1__8_ ( .D(n110), .CK(clk), .Q(queueRegister[18]) );
  DFFSHQX8TS queueEndPointer_reg_8_ ( .D(n424), .CK(clk), .SN(n447), .Q(n437)
         );
  DFFHQX4TS queueRegister_reg_6__8_ ( .D(n1050), .CK(clk), .Q(
        queueRegister[68]) );
  DFFHQX4TS queueRegister_reg_6__7_ ( .D(n112), .CK(clk), .Q(queueRegister[67]) );
  DFFHQX4TS queueRegister_reg_6__5_ ( .D(n1260), .CK(clk), .Q(
        queueRegister[65]) );
  DFFHQX4TS queueRegister_reg_6__2_ ( .D(n147), .CK(clk), .Q(queueRegister[62]) );
  DFFHQX4TS queueRegister_reg_6__1_ ( .D(n154), .CK(clk), .Q(queueRegister[61]) );
  DFFHQX4TS queueRegister_reg_0__8_ ( .D(n111), .CK(clk), .Q(queueRegister[8])
         );
  DFFSHQX8TS queueEndPointer_reg_5_ ( .D(n426), .CK(clk), .SN(n447), .Q(n433)
         );
  DFFRX4TS queueEndPointer_reg_2_ ( .D(n181), .CK(clk), .RN(n447), .Q(
        queueEndPointer[2]), .QN(n435) );
  DFFRHQX2TS queueRegister_reg_4__0_ ( .D(n163), .CK(clk), .RN(1'b1), .Q(
        queueRegister[40]) );
  DFFRHQX2TS queueRegister_reg_1__0_ ( .D(n166), .CK(clk), .RN(1'b1), .Q(
        queueRegister[10]) );
  DFFSX4TS queueEndPointer_reg_0_ ( .D(n195), .CK(clk), .SN(n447), .Q(n430) );
  DFFHQX4TS queueRegister_reg_3__9_ ( .D(n171), .CK(clk), .Q(queueRegister[39]) );
  DFFHQX4TS queueRegister_reg_3__4_ ( .D(n136), .CK(clk), .Q(queueRegister[34]) );
  DFFHQX4TS queueRegister_reg_3__2_ ( .D(n150), .CK(clk), .Q(queueRegister[32]) );
  DFFHQX4TS queueRegister_reg_6__9_ ( .D(n168), .CK(clk), .Q(queueRegister[69]) );
  DFFHQX4TS queueRegister_reg_5__9_ ( .D(n169), .CK(clk), .Q(queueRegister[59]) );
  DFFHQX4TS queueRegister_reg_5__2_ ( .D(n148), .CK(clk), .Q(queueRegister[52]) );
  DFFNSRX1TS queueFrontPointerBuffer_reg_1_ ( .D(n93), .CKN(n210), .SN(1'b1), 
        .RN(n83), .Q(queueFrontPointerBuffer[1]), .QN(n408) );
  DFFHQX4TS queueRegister_reg_6__4_ ( .D(n404), .CK(clk), .Q(queueRegister[64]) );
  DFFHQX4TS queueRegister_reg_0__0_ ( .D(n403), .CK(clk), .Q(queueRegister[0])
         );
  DFFQX2TS queueRegister_reg_2__1_ ( .D(n158), .CK(clk), .Q(queueRegister[21])
         );
  TLATX4TS finished_reg ( .G(N89), .D(N90), .Q(finished), .QN(n409) );
  DFFSHQX1TS queueEndPointer_reg_6_ ( .D(n427), .CK(clk), .SN(n447), .Q(n432)
         );
  DFFSHQX1TS queueEndPointer_reg_4_ ( .D(n405), .CK(clk), .SN(n447), .Q(n411)
         );
  MX2X1TS U201 ( .A(n361), .B(queueRegister[53]), .S0(n387), .Y(n141) );
  NOR2BX1TS U202 ( .AN(n254), .B(n194), .Y(n214) );
  CLKINVX2TS U203 ( .A(n244), .Y(n363) );
  NAND2X6TS U204 ( .A(n268), .B(n241), .Y(n388) );
  CLKINVX2TS U205 ( .A(n280), .Y(n261) );
  NOR2BX2TS U206 ( .AN(n444), .B(finished), .Y(n375) );
  CLKINVX2TS U207 ( .A(n273), .Y(n272) );
  NOR2X1TS U208 ( .A(n446), .B(n435), .Y(n227) );
  NAND2X1TS U209 ( .A(queueEndPointer[5]), .B(queueEndPointer[4]), .Y(n347) );
  INVX2TS U210 ( .A(n437), .Y(queueEndPointer[8]) );
  INVX2TS U211 ( .A(n433), .Y(queueEndPointer[5]) );
  BUFX4TS U212 ( .A(indexCounter[5]), .Y(n364) );
  AND2X2TS U213 ( .A(n432), .B(n197), .Y(n234) );
  CLKBUFX2TS U214 ( .A(resetInputQueue), .Y(n298) );
  MX2X1TS U215 ( .A(n361), .B(queueRegister[43]), .S0(n390), .Y(n142) );
  MX2X1TS U216 ( .A(n361), .B(queueRegister[13]), .S0(n386), .Y(n145) );
  MX2X1TS U217 ( .A(n361), .B(queueRegister[3]), .S0(n389), .Y(n146) );
  MX2X1TS U218 ( .A(n361), .B(queueRegister[23]), .S0(n388), .Y(n144) );
  MX2X1TS U219 ( .A(n361), .B(queueRegister[63]), .S0(n383), .Y(n140) );
  MX2X1TS U220 ( .A(n361), .B(queueRegister[33]), .S0(n385), .Y(n143) );
  CLKINVX3TS U221 ( .A(n206), .Y(n343) );
  OAI21XLTS U222 ( .A0(n247), .A1(finished), .B0(n246), .Y(n1010) );
  NAND2X2TS U223 ( .A(n338), .B(n337), .Y(n357) );
  NAND3BX1TS U224 ( .AN(n347), .B(n343), .C(n342), .Y(n344) );
  NAND2X6TS U225 ( .A(n238), .B(n239), .Y(n226) );
  CLKINVX3TS U226 ( .A(n389), .Y(n201) );
  NAND2X8TS U227 ( .A(n200), .B(n199), .Y(n389) );
  NOR2X8TS U228 ( .A(n196), .B(n226), .Y(n200) );
  NOR2X8TS U229 ( .A(n226), .B(n225), .Y(n231) );
  NAND2X6TS U230 ( .A(n218), .B(n236), .Y(n225) );
  NAND2BX4TS U231 ( .AN(finished), .B(pixelValue), .Y(n367) );
  BUFX6TS U232 ( .A(indexCounter[8]), .Y(n365) );
  NOR2X4TS U233 ( .A(n241), .B(n435), .Y(n219) );
  CLKINVX12TS U234 ( .A(n240), .Y(n268) );
  XNOR2X1TS U235 ( .A(n186), .B(n361), .Y(n247) );
  NOR2BX2TS U236 ( .AN(n363), .B(n280), .Y(n186) );
  NAND2BX2TS U237 ( .AN(n269), .B(queueRegister[30]), .Y(n270) );
  CLKINVX1TS U238 ( .A(n385), .Y(n269) );
  AND2X8TS U239 ( .A(n235), .B(n234), .Y(n237) );
  OAI21X1TS U240 ( .A0(n279), .A1(finished), .B0(n278), .Y(n97) );
  NAND2X2TS U241 ( .A(queueEndPointer[6]), .B(queueEndPointer[7]), .Y(n336) );
  OAI2BB1X2TS U242 ( .A0N(n386), .A1N(queueRegister[10]), .B0(n233), .Y(n166)
         );
  OAI2BB1X2TS U243 ( .A0N(n390), .A1N(queueRegister[40]), .B0(n229), .Y(n163)
         );
  NAND3X4TS U244 ( .A(n211), .B(indexCounter[0]), .C(n372), .Y(n273) );
  AND4X2TS U245 ( .A(n384), .B(n372), .C(indexCounter[0]), .D(n371), .Y(n376)
         );
  NAND2X4TS U246 ( .A(n372), .B(indexCounter[0]), .Y(n280) );
  INVX1TS U247 ( .A(n214), .Y(n215) );
  AND2X4TS U248 ( .A(n434), .B(n411), .Y(n238) );
  OR2X1TS U249 ( .A(queueEndPointer[8]), .B(n369), .Y(n339) );
  INVX2TS U250 ( .A(n245), .Y(n246) );
  XOR2X1TS U251 ( .A(n435), .B(n342), .Y(n185) );
  CLKINVX3TS U252 ( .A(n192), .Y(n193) );
  MX2X2TS U253 ( .A(queueRegister[64]), .B(n391), .S0(n223), .Y(n404) );
  NAND2X6TS U254 ( .A(n231), .B(n230), .Y(n386) );
  NAND2X6TS U255 ( .A(n231), .B(n227), .Y(n390) );
  INVX1TS U256 ( .A(n388), .Y(n242) );
  NAND2X6TS U257 ( .A(n205), .B(n204), .Y(n383) );
  CLKINVX2TS U258 ( .A(n265), .Y(n266) );
  INVX1TS U259 ( .A(n249), .Y(n250) );
  XOR2X1TS U260 ( .A(n344), .B(n432), .Y(n346) );
  CLKINVX2TS U261 ( .A(n442), .Y(n263) );
  CLKBUFX2TS U262 ( .A(dequeue), .Y(n210) );
  INVX3TS U263 ( .A(n225), .Y(n220) );
  MX2X2TS U264 ( .A(n365), .B(queueRegister[8]), .S0(n389), .Y(n111) );
  INVX1TS U265 ( .A(n209), .Y(n405) );
  NAND2BX1TS U266 ( .AN(n369), .B(n433), .Y(n355) );
  INVX2TS U267 ( .A(n409), .Y(n254) );
  OR2X2TS U268 ( .A(n445), .B(n409), .Y(n278) );
  NOR2X2TS U269 ( .A(n357), .B(n437), .Y(n358) );
  OR2X4TS U270 ( .A(n376), .B(n444), .Y(n382) );
  NAND2X4TS U271 ( .A(n342), .B(n343), .Y(n353) );
  INVX1TS U272 ( .A(n347), .Y(n348) );
  NAND2X6TS U273 ( .A(n364), .B(n391), .Y(n274) );
  CLKINVX2TS U274 ( .A(n432), .Y(queueEndPointer[6]) );
  CLKINVX2TS U275 ( .A(n413), .Y(n189) );
  CLKBUFX2TS U276 ( .A(n384), .Y(n188) );
  NAND2X4TS U277 ( .A(n446), .B(queueEndPointer[1]), .Y(n282) );
  NOR2X4TS U278 ( .A(n273), .B(n414), .Y(n248) );
  NAND2X2TS U279 ( .A(n341), .B(n228), .Y(n229) );
  NAND2X2TS U280 ( .A(n341), .B(n232), .Y(n233) );
  CLKINVX1TS U281 ( .A(n341), .Y(n187) );
  INVX3TS U282 ( .A(n211), .Y(n192) );
  CLKINVX6TS U283 ( .A(n439), .Y(n361) );
  OAI21XLTS U284 ( .A0(n258), .A1(finished), .B0(n257), .Y(n1030) );
  XOR2X4TS U285 ( .A(n248), .B(n443), .Y(n251) );
  CLKINVX6TS U286 ( .A(n274), .Y(n373) );
  NAND4X4TS U287 ( .A(n220), .B(n239), .C(n238), .D(n219), .Y(n387) );
  BUFX6TS U288 ( .A(indexCounter[1]), .Y(n372) );
  CLKINVX6TS U289 ( .A(n440), .Y(n341) );
  INVX2TS U290 ( .A(n383), .Y(n223) );
  MX2X1TS U291 ( .A(queueRegister[0]), .B(indexCounter[0]), .S0(n201), .Y(n403) );
  INVX2TS U292 ( .A(n386), .Y(n232) );
  INVX2TS U293 ( .A(n390), .Y(n228) );
  MX2X1TS U294 ( .A(n372), .B(queueRegister[61]), .S0(n383), .Y(n154) );
  MX2X1TS U295 ( .A(n363), .B(queueRegister[62]), .S0(n383), .Y(n147) );
  MX2X1TS U296 ( .A(n364), .B(queueRegister[65]), .S0(n383), .Y(n1260) );
  MX2X1TS U297 ( .A(n371), .B(queueRegister[67]), .S0(n383), .Y(n112) );
  MX2X1TS U298 ( .A(n365), .B(queueRegister[68]), .S0(n383), .Y(n1050) );
  MX2X1TS U299 ( .A(n365), .B(queueRegister[18]), .S0(n386), .Y(n110) );
  MX2X1TS U300 ( .A(n371), .B(queueRegister[17]), .S0(n386), .Y(n117) );
  MX2X1TS U301 ( .A(n364), .B(queueRegister[45]), .S0(n390), .Y(n128) );
  MX2X1TS U302 ( .A(n372), .B(queueRegister[11]), .S0(n386), .Y(n159) );
  MX2X1TS U303 ( .A(indexCounter[9]), .B(queueRegister[49]), .S0(n390), .Y(
        n170) );
  MX2X1TS U304 ( .A(n363), .B(queueRegister[42]), .S0(n390), .Y(n149) );
  MX2X1TS U305 ( .A(n371), .B(queueRegister[47]), .S0(n390), .Y(n114) );
  MX2X1TS U306 ( .A(n365), .B(queueRegister[48]), .S0(n390), .Y(n1070) );
  MX2X1TS U307 ( .A(n391), .B(queueRegister[14]), .S0(n386), .Y(n138) );
  MX2X1TS U308 ( .A(n384), .B(queueRegister[16]), .S0(n386), .Y(n124) );
  MX2X1TS U309 ( .A(n391), .B(queueRegister[44]), .S0(n390), .Y(n135) );
  MX2X1TS U310 ( .A(n384), .B(queueRegister[46]), .S0(n390), .Y(n121) );
  MX2X1TS U311 ( .A(indexCounter[9]), .B(queueRegister[19]), .S0(n386), .Y(
        n173) );
  MX2X1TS U312 ( .A(n364), .B(queueRegister[15]), .S0(n386), .Y(n131) );
  MX2X1TS U313 ( .A(n372), .B(queueRegister[41]), .S0(n390), .Y(n156) );
  INVX2TS U314 ( .A(n387), .Y(n221) );
  MX2X1TS U315 ( .A(n362), .B(queueRegister[22]), .S0(n388), .Y(n151) );
  MX2X1TS U316 ( .A(n362), .B(queueRegister[12]), .S0(n386), .Y(n152) );
  MX2X1TS U317 ( .A(n365), .B(queueRegister[58]), .S0(n387), .Y(n1060) );
  MX2X1TS U318 ( .A(n371), .B(queueRegister[57]), .S0(n387), .Y(n113) );
  MX2X1TS U319 ( .A(n372), .B(queueRegister[51]), .S0(n387), .Y(n155) );
  MX2X1TS U320 ( .A(n364), .B(queueRegister[55]), .S0(n387), .Y(n1270) );
  MX2X1TS U321 ( .A(n362), .B(queueRegister[52]), .S0(n387), .Y(n148) );
  MX2X1TS U322 ( .A(indexCounter[9]), .B(queueRegister[59]), .S0(n387), .Y(
        n169) );
  MX2X1TS U323 ( .A(n384), .B(queueRegister[56]), .S0(n387), .Y(n120) );
  MX2X1TS U324 ( .A(n391), .B(queueRegister[54]), .S0(n387), .Y(n134) );
  MX2X1TS U325 ( .A(indexCounter[9]), .B(queueRegister[69]), .S0(n383), .Y(
        n168) );
  MX2X1TS U326 ( .A(n384), .B(queueRegister[66]), .S0(n383), .Y(n119) );
  MX2X1TS U327 ( .A(n189), .B(queueRegister[31]), .S0(n385), .Y(n157) );
  MX2X1TS U328 ( .A(n362), .B(queueRegister[32]), .S0(n385), .Y(n150) );
  MX2X1TS U329 ( .A(n365), .B(queueRegister[38]), .S0(n385), .Y(n108) );
  MX2X1TS U330 ( .A(n371), .B(queueRegister[37]), .S0(n385), .Y(n115) );
  MX2X1TS U331 ( .A(n364), .B(queueRegister[35]), .S0(n385), .Y(n129) );
  MX2X1TS U332 ( .A(n384), .B(queueRegister[36]), .S0(n385), .Y(n122) );
  MX2X1TS U333 ( .A(n391), .B(queueRegister[34]), .S0(n385), .Y(n136) );
  MX2X1TS U334 ( .A(indexCounter[9]), .B(queueRegister[39]), .S0(n385), .Y(
        n171) );
  MX2X1TS U335 ( .A(n365), .B(queueRegister[28]), .S0(n388), .Y(n109) );
  MX2X1TS U336 ( .A(n371), .B(queueRegister[27]), .S0(n388), .Y(n116) );
  MX2X1TS U337 ( .A(n372), .B(queueRegister[21]), .S0(n388), .Y(n158) );
  MX2X1TS U338 ( .A(n371), .B(queueRegister[7]), .S0(n389), .Y(n118) );
  MX2X1TS U339 ( .A(n372), .B(queueRegister[1]), .S0(n389), .Y(n160) );
  MX2X1TS U340 ( .A(n364), .B(queueRegister[25]), .S0(n388), .Y(n130) );
  MX2X1TS U341 ( .A(indexCounter[9]), .B(queueRegister[29]), .S0(n388), .Y(
        n172) );
  MX2X1TS U342 ( .A(n364), .B(queueRegister[5]), .S0(n389), .Y(n132) );
  MX2X1TS U343 ( .A(n363), .B(queueRegister[2]), .S0(n389), .Y(n153) );
  MX2X1TS U344 ( .A(indexCounter[9]), .B(queueRegister[9]), .S0(n389), .Y(n174) );
  MX2X1TS U345 ( .A(n384), .B(queueRegister[26]), .S0(n388), .Y(n123) );
  MX2X1TS U346 ( .A(n391), .B(queueRegister[4]), .S0(n389), .Y(n139) );
  INVX1TS U347 ( .A(n256), .Y(n257) );
  XNOR2X1TS U348 ( .A(n341), .B(n189), .Y(n258) );
  NOR2BX1TS U349 ( .AN(finished), .B(n413), .Y(n256) );
  OAI21XLTS U350 ( .A0(n255), .A1(n254), .B0(n253), .Y(n1000) );
  INVX1TS U351 ( .A(n252), .Y(n253) );
  NOR2BX1TS U352 ( .AN(n254), .B(n414), .Y(n252) );
  NOR2BX1TS U353 ( .AN(finished), .B(n443), .Y(n249) );
  CLKINVX1TS U354 ( .A(n362), .Y(n190) );
  CLKINVX3TS U355 ( .A(n441), .Y(n362) );
  CLKINVX1TS U356 ( .A(indexCounter[2]), .Y(n244) );
  INVX2TS U357 ( .A(n192), .Y(n191) );
  NOR2BX1TS U358 ( .AN(finished), .B(n439), .Y(n245) );
  XOR2X1TS U359 ( .A(n273), .B(n391), .Y(n255) );
  NOR2X4TS U360 ( .A(n273), .B(n274), .Y(n213) );
  INVX2TS U361 ( .A(n367), .Y(n369) );
  XNOR2X1TS U362 ( .A(n446), .B(n369), .Y(n195) );
  INVX2TS U363 ( .A(n411), .Y(queueEndPointer[4]) );
  INVX2TS U364 ( .A(n298), .Y(n447) );
  NOR2X8TS U365 ( .A(queueEndPointer[7]), .B(queueEndPointer[5]), .Y(n236) );
  INVX2TS U366 ( .A(n236), .Y(n196) );
  NOR2X8TS U367 ( .A(queueEndPointer[8]), .B(queueEndPointer[9]), .Y(n239) );
  INVX8TS U368 ( .A(n430), .Y(n446) );
  OR2X4TS U369 ( .A(n446), .B(queueEndPointer[2]), .Y(n198) );
  NOR2X1TS U370 ( .A(n367), .B(n298), .Y(n197) );
  NAND2X2TS U371 ( .A(n234), .B(n436), .Y(n217) );
  NOR2X2TS U372 ( .A(n198), .B(n217), .Y(n199) );
  BUFX6TS U373 ( .A(indexCounter[4]), .Y(n391) );
  INVX2TS U374 ( .A(n234), .Y(n202) );
  NAND3BX4TS U375 ( .AN(n202), .B(n238), .C(n236), .Y(n203) );
  NOR2BX4TS U376 ( .AN(n239), .B(n203), .Y(n205) );
  NOR3X2TS U377 ( .A(n446), .B(n435), .C(n436), .Y(n204) );
  CLKINVX6TS U378 ( .A(n282), .Y(n342) );
  NAND2X2TS U379 ( .A(queueEndPointer[3]), .B(queueEndPointer[2]), .Y(n206) );
  CLKINVX6TS U380 ( .A(n353), .Y(n337) );
  XOR2X1TS U381 ( .A(n337), .B(n411), .Y(n208) );
  NAND2X1TS U382 ( .A(queueEndPointer[4]), .B(n367), .Y(n207) );
  OAI21X1TS U383 ( .A0(n208), .A1(n367), .B0(n207), .Y(n209) );
  BUFX6TS U386 ( .A(writeBufferEnable), .Y(n429) );
  NAND2X2TS U387 ( .A(indexCounter[2]), .B(indexCounter[3]), .Y(n260) );
  CLKINVX6TS U388 ( .A(n260), .Y(n211) );
  INVX2TS U389 ( .A(indexCounter[6]), .Y(n212) );
  CLKINVX6TS U390 ( .A(n212), .Y(n384) );
  XNOR2X4TS U391 ( .A(n213), .B(n188), .Y(n216) );
  OAI21X2TS U392 ( .A0(n216), .A1(n254), .B0(n215), .Y(n980) );
  INVX2TS U393 ( .A(n217), .Y(n218) );
  INVX4TS U394 ( .A(n446), .Y(n241) );
  NAND2X1TS U395 ( .A(n341), .B(n221), .Y(n222) );
  OAI2BB1X2TS U396 ( .A0N(n387), .A1N(queueRegister[50]), .B0(n222), .Y(n162)
         );
  NAND2X1TS U397 ( .A(n341), .B(n223), .Y(n224) );
  OAI2BB1X2TS U398 ( .A0N(n383), .A1N(queueRegister[60]), .B0(n224), .Y(n161)
         );
  NOR2X2TS U399 ( .A(queueEndPointer[2]), .B(n241), .Y(n230) );
  NOR2X4TS U400 ( .A(queueEndPointer[2]), .B(n436), .Y(n235) );
  NAND4X4TS U401 ( .A(n239), .B(n238), .C(n237), .D(n236), .Y(n240) );
  NAND2X1TS U402 ( .A(n341), .B(n242), .Y(n243) );
  OAI2BB1X2TS U403 ( .A0N(n388), .A1N(queueRegister[20]), .B0(n243), .Y(n165)
         );
  OAI21X2TS U404 ( .A0(n251), .A1(finished), .B0(n250), .Y(n990) );
  BUFX6TS U405 ( .A(indexCounter[7]), .Y(n371) );
  NAND3X4TS U406 ( .A(n365), .B(n371), .C(n384), .Y(n259) );
  INVX2TS U407 ( .A(n259), .Y(n262) );
  NAND4X4TS U408 ( .A(n262), .B(n261), .C(n373), .D(n193), .Y(n264) );
  XOR2X4TS U409 ( .A(n264), .B(n263), .Y(n267) );
  NOR2BX1TS U410 ( .AN(finished), .B(n442), .Y(n265) );
  OAI21X2TS U411 ( .A0(n267), .A1(finished), .B0(n266), .Y(n95) );
  NAND2X6TS U412 ( .A(n268), .B(n446), .Y(n385) );
  OAI21X1TS U413 ( .A0(n385), .A1(n440), .B0(n270), .Y(n164) );
  AND2X2TS U414 ( .A(n371), .B(n384), .Y(n271) );
  NAND3X2TS U415 ( .A(n272), .B(n373), .C(n271), .Y(n277) );
  OAI21X1TS U416 ( .A0(n194), .A1(n273), .B0(n445), .Y(n276) );
  NAND2X1TS U417 ( .A(n274), .B(n445), .Y(n275) );
  NAND3X2TS U418 ( .A(n277), .B(n276), .C(n275), .Y(n279) );
  XOR2X1TS U419 ( .A(n362), .B(n280), .Y(n281) );
  MXI2X1TS U420 ( .A(n281), .B(n190), .S0(finished), .Y(n1020) );
  MXI2X1TS U421 ( .A(n185), .B(n435), .S0(n367), .Y(n181) );
  INVX1TS U422 ( .A(resetBuffer), .Y(n81) );
  NOR2X2TS U423 ( .A(queueFrontPointerBuffer[2]), .B(n408), .Y(n332) );
  NOR2X2TS U424 ( .A(queueFrontPointerBuffer[2]), .B(
        queueFrontPointerBuffer[1]), .Y(n331) );
  NOR2X1TS U425 ( .A(queueFrontPointerBuffer[1]), .B(n415), .Y(n330) );
  AOI222XLTS U426 ( .A0(n332), .A1(queueRegisterBuffer[35]), .B0(n331), .B1(
        queueRegisterBuffer[15]), .C0(n330), .C1(queueRegisterBuffer[55]), .Y(
        n285) );
  NOR2X1TS U427 ( .A(n415), .B(n408), .Y(n394) );
  AOI222XLTS U428 ( .A0(n332), .A1(queueRegisterBuffer[25]), .B0(n331), .B1(
        queueRegisterBuffer[5]), .C0(n330), .C1(queueRegisterBuffer[45]), .Y(
        n283) );
  AOI2BB2XLTS U429 ( .B0(n394), .B1(queueRegisterBuffer[65]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n283), .Y(n284) );
  OAI21XLTS U430 ( .A0(n285), .A1(n423), .B0(n284), .Y(N102) );
  AOI222XLTS U431 ( .A0(n332), .A1(queueRegisterBuffer[34]), .B0(n331), .B1(
        queueRegisterBuffer[14]), .C0(n330), .C1(queueRegisterBuffer[54]), .Y(
        n288) );
  AOI222XLTS U432 ( .A0(n332), .A1(queueRegisterBuffer[24]), .B0(n331), .B1(
        queueRegisterBuffer[4]), .C0(n330), .C1(queueRegisterBuffer[44]), .Y(
        n286) );
  AOI2BB2XLTS U433 ( .B0(n394), .B1(queueRegisterBuffer[64]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n286), .Y(n287) );
  OAI21XLTS U434 ( .A0(n288), .A1(n423), .B0(n287), .Y(N103) );
  AOI222XLTS U435 ( .A0(n332), .A1(queueRegisterBuffer[33]), .B0(n331), .B1(
        queueRegisterBuffer[13]), .C0(n330), .C1(queueRegisterBuffer[53]), .Y(
        n291) );
  AOI222XLTS U436 ( .A0(n332), .A1(queueRegisterBuffer[23]), .B0(n331), .B1(
        queueRegisterBuffer[3]), .C0(n330), .C1(queueRegisterBuffer[43]), .Y(
        n289) );
  AOI2BB2XLTS U437 ( .B0(n394), .B1(queueRegisterBuffer[63]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n289), .Y(n290) );
  OAI21XLTS U438 ( .A0(n291), .A1(n423), .B0(n290), .Y(N104) );
  AOI222XLTS U439 ( .A0(n332), .A1(queueRegisterBuffer[37]), .B0(n331), .B1(
        queueRegisterBuffer[17]), .C0(n330), .C1(queueRegisterBuffer[57]), .Y(
        n294) );
  AOI222XLTS U440 ( .A0(n332), .A1(queueRegisterBuffer[27]), .B0(n331), .B1(
        queueRegisterBuffer[7]), .C0(n330), .C1(queueRegisterBuffer[47]), .Y(
        n292) );
  AOI2BB2XLTS U441 ( .B0(n394), .B1(queueRegisterBuffer[67]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n292), .Y(n293) );
  OAI21XLTS U442 ( .A0(n294), .A1(n423), .B0(n293), .Y(N100) );
  AOI222XLTS U443 ( .A0(n332), .A1(queueRegisterBuffer[36]), .B0(n331), .B1(
        queueRegisterBuffer[16]), .C0(n330), .C1(queueRegisterBuffer[56]), .Y(
        n297) );
  AOI222XLTS U444 ( .A0(n332), .A1(queueRegisterBuffer[26]), .B0(n331), .B1(
        queueRegisterBuffer[6]), .C0(n330), .C1(queueRegisterBuffer[46]), .Y(
        n295) );
  AOI2BB2XLTS U445 ( .B0(n394), .B1(queueRegisterBuffer[66]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n295), .Y(n296) );
  OAI21XLTS U446 ( .A0(n297), .A1(n423), .B0(n296), .Y(N101) );
  NAND4XLTS U447 ( .A(n362), .B(n445), .C(n194), .D(n447), .Y(n301) );
  NOR4XLTS U448 ( .A(n364), .B(n391), .C(n361), .D(n365), .Y(n299) );
  NAND3XLTS U449 ( .A(n189), .B(n299), .C(n187), .Y(n300) );
  NOR3XLTS U450 ( .A(indexCounter[9]), .B(n301), .C(n300), .Y(N90) );
  AOI222XLTS U451 ( .A0(n332), .A1(queueRegisterBuffer[38]), .B0(n331), .B1(
        queueRegisterBuffer[18]), .C0(n330), .C1(queueRegisterBuffer[58]), .Y(
        n304) );
  AOI222XLTS U452 ( .A0(n332), .A1(queueRegisterBuffer[28]), .B0(n331), .B1(
        queueRegisterBuffer[8]), .C0(n330), .C1(queueRegisterBuffer[48]), .Y(
        n302) );
  AOI2BB2XLTS U453 ( .B0(n394), .B1(queueRegisterBuffer[68]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n302), .Y(n303) );
  OAI21XLTS U454 ( .A0(n304), .A1(n423), .B0(n303), .Y(N99) );
  AOI222XLTS U455 ( .A0(n332), .A1(queueRegisterBuffer[32]), .B0(n331), .B1(
        queueRegisterBuffer[12]), .C0(n330), .C1(queueRegisterBuffer[52]), .Y(
        n307) );
  AOI222XLTS U456 ( .A0(n332), .A1(queueRegisterBuffer[22]), .B0(n331), .B1(
        queueRegisterBuffer[2]), .C0(n330), .C1(queueRegisterBuffer[42]), .Y(
        n305) );
  AOI2BB2XLTS U457 ( .B0(n394), .B1(queueRegisterBuffer[62]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n305), .Y(n306) );
  OAI21XLTS U458 ( .A0(n307), .A1(n423), .B0(n306), .Y(N105) );
  AOI222XLTS U459 ( .A0(n332), .A1(queueRegisterBuffer[31]), .B0(n331), .B1(
        queueRegisterBuffer[11]), .C0(n330), .C1(queueRegisterBuffer[51]), .Y(
        n310) );
  AOI222XLTS U460 ( .A0(n332), .A1(queueRegisterBuffer[21]), .B0(n331), .B1(
        queueRegisterBuffer[1]), .C0(n330), .C1(queueRegisterBuffer[41]), .Y(
        n308) );
  AOI2BB2XLTS U461 ( .B0(n394), .B1(queueRegisterBuffer[61]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n308), .Y(n309) );
  OAI21XLTS U462 ( .A0(n310), .A1(n423), .B0(n309), .Y(N106) );
  AOI222XLTS U463 ( .A0(n332), .A1(queueRegisterBuffer[39]), .B0(n331), .B1(
        queueRegisterBuffer[19]), .C0(n330), .C1(queueRegisterBuffer[59]), .Y(
        n313) );
  AOI222XLTS U464 ( .A0(n332), .A1(queueRegisterBuffer[29]), .B0(n331), .B1(
        queueRegisterBuffer[9]), .C0(n330), .C1(queueRegisterBuffer[49]), .Y(
        n311) );
  AOI2BB2XLTS U465 ( .B0(n394), .B1(queueRegisterBuffer[69]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n311), .Y(n312) );
  OAI21XLTS U466 ( .A0(n313), .A1(n423), .B0(n312), .Y(N98) );
  XOR2XLTS U467 ( .A(n418), .B(queueEndPointerBuffer[3]), .Y(n315) );
  XOR2XLTS U468 ( .A(n415), .B(queueEndPointerBuffer[2]), .Y(n314) );
  NAND2X1TS U469 ( .A(n315), .B(n314), .Y(n329) );
  XOR2XLTS U470 ( .A(n417), .B(queueEndPointerBuffer[6]), .Y(n317) );
  XOR2XLTS U471 ( .A(n408), .B(queueEndPointerBuffer[1]), .Y(n316) );
  NAND2X1TS U472 ( .A(n317), .B(n316), .Y(n328) );
  XOR2XLTS U473 ( .A(n421), .B(queueEndPointerBuffer[8]), .Y(n319) );
  XOR2XLTS U474 ( .A(n422), .B(queueEndPointerBuffer[5]), .Y(n318) );
  NAND2X1TS U475 ( .A(n319), .B(n318), .Y(n327) );
  NOR2X1TS U476 ( .A(resetBuffer), .B(n429), .Y(n83) );
  XNOR2X1TS U477 ( .A(n423), .B(queueEndPointerBuffer[0]), .Y(n321) );
  XNOR2X1TS U478 ( .A(n419), .B(queueEndPointerBuffer[9]), .Y(n320) );
  NOR2XLTS U479 ( .A(n321), .B(n320), .Y(n325) );
  XNOR2X1TS U480 ( .A(n416), .B(queueEndPointerBuffer[4]), .Y(n323) );
  XNOR2X1TS U481 ( .A(n420), .B(queueEndPointerBuffer[7]), .Y(n322) );
  NOR2XLTS U482 ( .A(n323), .B(n322), .Y(n324) );
  NAND3XLTS U483 ( .A(n83), .B(n325), .C(n324), .Y(n326) );
  NOR4XLTS U484 ( .A(n329), .B(n328), .C(n327), .D(n326), .Y(N127) );
  AOI222XLTS U485 ( .A0(n332), .A1(queueRegisterBuffer[30]), .B0(n331), .B1(
        queueRegisterBuffer[10]), .C0(n330), .C1(queueRegisterBuffer[50]), .Y(
        n335) );
  AOI222XLTS U486 ( .A0(n332), .A1(queueRegisterBuffer[20]), .B0(n331), .B1(
        queueRegisterBuffer[0]), .C0(n330), .C1(queueRegisterBuffer[40]), .Y(
        n333) );
  AOI2BB2XLTS U487 ( .B0(n394), .B1(queueRegisterBuffer[60]), .A0N(
        queueFrontPointerBuffer[0]), .A1N(n333), .Y(n334) );
  OAI21XLTS U488 ( .A0(n335), .A1(n423), .B0(n334), .Y(N107) );
  NOR2X2TS U489 ( .A(n347), .B(n336), .Y(n338) );
  XOR2X1TS U490 ( .A(n357), .B(n437), .Y(n340) );
  OAI21X1TS U491 ( .A0(n340), .A1(n367), .B0(n339), .Y(n424) );
  XOR2X1TS U492 ( .A(n409), .B(n341), .Y(n1040) );
  NAND2BX1TS U493 ( .AN(n369), .B(n432), .Y(n345) );
  OAI21X1TS U494 ( .A0(n346), .A1(n367), .B0(n345), .Y(n427) );
  NAND2X1TS U495 ( .A(n348), .B(queueEndPointer[6]), .Y(n349) );
  NOR2X1TS U496 ( .A(n353), .B(n349), .Y(n350) );
  XNOR2X1TS U497 ( .A(n350), .B(n431), .Y(n352) );
  NAND2BX1TS U498 ( .AN(n369), .B(n431), .Y(n351) );
  OAI21X1TS U499 ( .A0(n352), .A1(n367), .B0(n351), .Y(n428) );
  NOR2X1TS U500 ( .A(n353), .B(n411), .Y(n354) );
  XNOR2X1TS U501 ( .A(n354), .B(n433), .Y(n356) );
  OAI21X1TS U502 ( .A0(n356), .A1(n367), .B0(n355), .Y(n426) );
  XNOR2X1TS U503 ( .A(n358), .B(n438), .Y(n360) );
  NAND2BX1TS U504 ( .AN(n369), .B(n438), .Y(n359) );
  OAI21X1TS U505 ( .A0(n360), .A1(n367), .B0(n359), .Y(n425) );
  NAND2BXLTS U506 ( .AN(N90), .B(n447), .Y(N89) );
  NAND2X1TS U507 ( .A(n342), .B(queueEndPointer[2]), .Y(n366) );
  XOR2X1TS U508 ( .A(n366), .B(n434), .Y(n368) );
  MXI2X1TS U509 ( .A(n368), .B(queueEndPointer[3]), .S0(n367), .Y(n410) );
  XOR2X1TS U510 ( .A(n436), .B(n446), .Y(n370) );
  CLKMX2X2TS U511 ( .A(n436), .B(n370), .S0(n369), .Y(n412) );
  NAND2X2TS U512 ( .A(n191), .B(n373), .Y(n379) );
  INVX2TS U513 ( .A(n379), .Y(n374) );
  NAND2X2TS U514 ( .A(n375), .B(n374), .Y(n377) );
  NAND2BX2TS U515 ( .AN(n377), .B(n376), .Y(n381) );
  NOR2X1TS U516 ( .A(n444), .B(n409), .Y(n378) );
  AOI21X2TS U517 ( .A0(n379), .A1(n365), .B0(n378), .Y(n380) );
  NAND3X1TS U518 ( .A(n382), .B(n381), .C(n380), .Y(n96) );
  CLKMX2X2TS U519 ( .A(n384), .B(queueRegister[6]), .S0(n389), .Y(n125) );
  CLKMX2X2TS U520 ( .A(n391), .B(queueRegister[24]), .S0(n388), .Y(n137) );
  NAND2BXLTS U521 ( .AN(N127), .B(n83), .Y(N126) );
  NOR2XLTS U522 ( .A(queueEmpty), .B(n423), .Y(n393) );
  AOI21X1TS U523 ( .A0(queueEmpty), .A1(n423), .B0(n393), .Y(n94) );
  AOI2BB2XLTS U524 ( .B0(queueFrontPointerBuffer[1]), .B1(n393), .A0N(n393), 
        .A1N(queueFrontPointerBuffer[1]), .Y(n93) );
  NAND2X1TS U525 ( .A(queueFrontPointerBuffer[1]), .B(n393), .Y(n392) );
  XNOR2X1TS U526 ( .A(queueFrontPointerBuffer[2]), .B(n392), .Y(n92) );
  NAND2X1TS U527 ( .A(n394), .B(n393), .Y(n396) );
  NAND3XLTS U528 ( .A(n394), .B(n393), .C(queueFrontPointerBuffer[3]), .Y(n397) );
  INVX2TS U529 ( .A(n397), .Y(n395) );
  AOI21X1TS U530 ( .A0(n396), .A1(n418), .B0(n395), .Y(n91) );
  NOR2XLTS U531 ( .A(n416), .B(n397), .Y(n398) );
  AOI21X1TS U532 ( .A0(n397), .A1(n416), .B0(n398), .Y(n900) );
  NAND2X1TS U533 ( .A(n398), .B(queueFrontPointerBuffer[5]), .Y(n399) );
  OA21XLTS U534 ( .A0(n398), .A1(queueFrontPointerBuffer[5]), .B0(n399), .Y(
        n890) );
  NOR2XLTS U535 ( .A(n417), .B(n399), .Y(n400) );
  AOI21X1TS U536 ( .A0(n399), .A1(n417), .B0(n400), .Y(n88) );
  NAND2X1TS U537 ( .A(n400), .B(queueFrontPointerBuffer[7]), .Y(n401) );
  OA21XLTS U538 ( .A0(n400), .A1(queueFrontPointerBuffer[7]), .B0(n401), .Y(
        n87) );
  XNOR2X1TS U539 ( .A(queueFrontPointerBuffer[8]), .B(n401), .Y(n86) );
  NAND2BXLTS U541 ( .AN(n401), .B(queueFrontPointerBuffer[8]), .Y(n402) );
  XNOR2X1TS U542 ( .A(queueFrontPointerBuffer[9]), .B(n402), .Y(n85) );
endmodule

