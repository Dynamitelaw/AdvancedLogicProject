
module softMax ( sumIn, result );
  input [99:0] sumIn;
  output [3:0] result;
  wire   n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;

  INVX2TS U605 ( .A(n881), .Y(n758) );
  NAND2BXLTS U606 ( .AN(n822), .B(n879), .Y(n831) );
  NAND2BXLTS U607 ( .AN(n1038), .B(n1110), .Y(n1044) );
  NAND2BXLTS U608 ( .AN(sumIn[24]), .B(n796), .Y(n801) );
  MXI2XLTS U609 ( .A(n1161), .B(n1160), .S0(n1286), .Y(n1219) );
  MXI2XLTS U610 ( .A(n1156), .B(n1155), .S0(n1180), .Y(n1222) );
  INVX2TS U611 ( .A(n1154), .Y(n1155) );
  MXI2XLTS U612 ( .A(n1151), .B(n1150), .S0(n1292), .Y(n1213) );
  INVX2TS U613 ( .A(n1149), .Y(n1150) );
  MXI2XLTS U614 ( .A(n1159), .B(n1158), .S0(n1292), .Y(n1223) );
  INVX2TS U615 ( .A(n1157), .Y(n1158) );
  INVX2TS U616 ( .A(n1222), .Y(n1224) );
  MXI2XLTS U617 ( .A(n1217), .B(n1216), .S0(n1232), .Y(n1218) );
  MXI2XLTS U618 ( .A(n1153), .B(n1152), .S0(n1285), .Y(n1221) );
  INVX2TS U619 ( .A(n1227), .Y(n676) );
  INVX2TS U620 ( .A(n1212), .Y(n677) );
  XOR2XLTS U621 ( .A(n664), .B(n663), .Y(n1234) );
  NAND2BXLTS U622 ( .AN(n751), .B(n886), .Y(n757) );
  AOI2BB1XLTS U623 ( .A0N(n839), .A1N(n864), .B0(n868), .Y(n807) );
  INVX2TS U624 ( .A(n882), .Y(n830) );
  XOR2XLTS U625 ( .A(n1032), .B(n1031), .Y(n1098) );
  OAI31X1TS U626 ( .A0(n960), .A1(n950), .A2(n952), .B0(n985), .Y(n943) );
  MXI2XLTS U627 ( .A(n1110), .B(n1109), .S0(n1108), .Y(n1152) );
  NAND2BXLTS U628 ( .AN(sumIn[84]), .B(n1009), .Y(n1014) );
  OAI31X1TS U629 ( .A0(n1027), .A1(n1026), .A2(n1025), .B0(n1024), .Y(n1090)
         );
  XOR2XLTS U630 ( .A(sumIn[83]), .B(n1021), .Y(n1092) );
  OAI31X1TS U631 ( .A0(n1030), .A1(n1037), .A2(n1028), .B0(n1065), .Y(n1021)
         );
  INVX2TS U632 ( .A(n1104), .Y(n1045) );
  XOR2XLTS U633 ( .A(n964), .B(n963), .Y(n1107) );
  XOR2XLTS U634 ( .A(n960), .B(n959), .Y(n1106) );
  NAND2BXLTS U635 ( .AN(n957), .B(n1103), .Y(n967) );
  OAI31X1TS U636 ( .A0(n949), .A1(n948), .A2(n947), .B0(n946), .Y(n1114) );
  INVX2TS U637 ( .A(n1113), .Y(n968) );
  XOR2XLTS U638 ( .A(n954), .B(n953), .Y(n1097) );
  OAI31X1TS U639 ( .A0(n941), .A1(n940), .A2(n945), .B0(n939), .Y(n1089) );
  NAND2BXLTS U640 ( .AN(sumIn[64]), .B(n932), .Y(n937) );
  OAI31X1TS U641 ( .A0(n740), .A1(n739), .A2(n737), .B0(n738), .Y(n869) );
  XOR2XLTS U642 ( .A(sumIn[43]), .B(n735), .Y(n871) );
  OAI31X1TS U643 ( .A0(n744), .A1(n750), .A2(n742), .B0(n741), .Y(n735) );
  OAI31X1TS U644 ( .A0(n813), .A1(n812), .A2(n810), .B0(n811), .Y(n889) );
  XOR2XLTS U645 ( .A(sumIn[23]), .B(n808), .Y(n891) );
  OAI31X1TS U646 ( .A0(n824), .A1(n815), .A2(n817), .B0(n814), .Y(n808) );
  XOR2XLTS U647 ( .A(n819), .B(n818), .Y(n873) );
  XOR2XLTS U648 ( .A(n828), .B(n827), .Y(n882) );
  XOR2XLTS U649 ( .A(n824), .B(n823), .Y(n883) );
  MXI2XLTS U650 ( .A(n886), .B(n885), .S0(n884), .Y(n1161) );
  XOR2XLTS U651 ( .A(n746), .B(n745), .Y(n875) );
  OAI31X1TS U652 ( .A0(n733), .A1(n732), .A2(n737), .B0(n731), .Y(n867) );
  NAND2BXLTS U653 ( .AN(sumIn[44]), .B(n723), .Y(n728) );
  INVX2TS U654 ( .A(n1174), .Y(n1175) );
  MXI2XLTS U655 ( .A(n1166), .B(n1165), .S0(n1164), .Y(n1215) );
  INVX2TS U656 ( .A(n1163), .Y(n1165) );
  INVX2TS U657 ( .A(n1213), .Y(n1214) );
  MXI2XLTS U658 ( .A(n1234), .B(n1233), .S0(n1232), .Y(n1235) );
  INVX2TS U659 ( .A(n1231), .Y(n1233) );
  AOI2BB1XLTS U660 ( .A0N(n1294), .A1N(n1221), .B0(n1220), .Y(n1230) );
  MXI2XLTS U661 ( .A(n1227), .B(n1226), .S0(n1246), .Y(n1228) );
  MXI2XLTS U662 ( .A(n1224), .B(n1223), .S0(n1199), .Y(n1229) );
  MXI2XLTS U663 ( .A(n1148), .B(n1147), .S0(n1164), .Y(n1210) );
  MXI2XLTS U664 ( .A(n1170), .B(n1169), .S0(n1285), .Y(n1208) );
  INVX2TS U665 ( .A(n1168), .Y(n1169) );
  OAI31X1TS U666 ( .A0(n662), .A1(n668), .A2(n660), .B0(n659), .Y(n653) );
  OAI31X1TS U667 ( .A0(n658), .A1(n657), .A2(n656), .B0(n655), .Y(n1211) );
  OAI31X1TS U668 ( .A0(n650), .A1(n649), .A2(n695), .B0(n648), .Y(n1244) );
  NAND2BXLTS U669 ( .AN(sumIn[4]), .B(n641), .Y(n646) );
  NAND2BXLTS U670 ( .AN(n669), .B(n1216), .Y(n675) );
  NAND2BXLTS U671 ( .AN(sumIn[56]), .B(n720), .Y(n708) );
  NAND2BXLTS U672 ( .AN(sumIn[46]), .B(n716), .Y(n706) );
  AOI2BB1XLTS U673 ( .A0N(n766), .A1N(n866), .B0(n867), .Y(n734) );
  MXI2XLTS U674 ( .A(n1089), .B(n1088), .S0(n1095), .Y(n1173) );
  INVX2TS U675 ( .A(n1054), .Y(n1083) );
  OAI31X1TS U676 ( .A0(n1018), .A1(n1017), .A2(n1023), .B0(n1016), .Y(n1087)
         );
  MXI2XLTS U677 ( .A(n1100), .B(n1099), .S0(n1284), .Y(n1149) );
  INVX2TS U678 ( .A(n1098), .Y(n1100) );
  MXI2XLTS U679 ( .A(n1093), .B(n1092), .S0(n1091), .Y(n1168) );
  INVX2TS U680 ( .A(n1090), .Y(n1093) );
  MXI2XLTS U681 ( .A(n1114), .B(n1113), .S0(n1283), .Y(n1170) );
  MXI2XLTS U682 ( .A(n1107), .B(n1106), .S0(n1283), .Y(n1159) );
  MXI2XLTS U683 ( .A(n1105), .B(n1104), .S0(n1284), .Y(n1157) );
  MXI2XLTS U684 ( .A(n1103), .B(n1102), .S0(n1101), .Y(n1153) );
  MXI2XLTS U685 ( .A(n1097), .B(n1096), .S0(n1095), .Y(n1151) );
  INVX2TS U686 ( .A(n1094), .Y(n1096) );
  NAND2BXLTS U687 ( .AN(sumIn[96]), .B(n1007), .Y(n1061) );
  NAND2BXLTS U688 ( .AN(sumIn[86]), .B(n1004), .Y(n1002) );
  XOR2XLTS U689 ( .A(n1005), .B(sumIn[86]), .Y(n1082) );
  INVX2TS U690 ( .A(n1107), .Y(n966) );
  AOI2BB1XLTS U691 ( .A0N(n976), .A1N(n1084), .B0(n1089), .Y(n942) );
  NAND2BXLTS U692 ( .AN(sumIn[76]), .B(n930), .Y(n982) );
  NAND2BXLTS U693 ( .AN(sumIn[66]), .B(n927), .Y(n925) );
  MXI2XLTS U694 ( .A(n864), .B(n863), .S0(n862), .Y(n1138) );
  MXI2XLTS U695 ( .A(n871), .B(n870), .S0(n1288), .Y(n1148) );
  INVX2TS U696 ( .A(n869), .Y(n870) );
  MXI2XLTS U697 ( .A(n891), .B(n890), .S0(n1287), .Y(n1147) );
  INVX2TS U698 ( .A(n889), .Y(n890) );
  MXI2XLTS U699 ( .A(n874), .B(n873), .S0(n900), .Y(n1163) );
  INVX2TS U700 ( .A(n872), .Y(n874) );
  MXI2XLTS U701 ( .A(n881), .B(n880), .S0(n1288), .Y(n1156) );
  MXI2XLTS U702 ( .A(n883), .B(n882), .S0(n900), .Y(n1154) );
  MXI2XLTS U703 ( .A(n879), .B(n878), .S0(n1287), .Y(n1160) );
  MXI2XLTS U704 ( .A(n877), .B(n876), .S0(n884), .Y(n1166) );
  INVX2TS U705 ( .A(n875), .Y(n876) );
  OAI31X1TS U706 ( .A0(n806), .A1(n805), .A2(n810), .B0(n804), .Y(n868) );
  MXI2XLTS U707 ( .A(n724), .B(n867), .S0(n884), .Y(n1146) );
  XOR2XLTS U708 ( .A(n790), .B(sumIn[26]), .Y(n902) );
  NAND2BXLTS U709 ( .AN(sumIn[36]), .B(n793), .Y(n781) );
  NAND2BXLTS U710 ( .AN(sumIn[26]), .B(n789), .Y(n779) );
  AO22XLTS U711 ( .A0(n1207), .A1(n1178), .B0(n1177), .B1(n1176), .Y(n1179) );
  AO21XLTS U712 ( .A0(n1177), .A1(n1175), .B0(n1176), .Y(n1178) );
  MXI2XLTS U713 ( .A(n1139), .B(n1138), .S0(n1180), .Y(n1204) );
  MXI2XLTS U714 ( .A(n1143), .B(n1142), .S0(n1141), .Y(n1202) );
  INVX2TS U715 ( .A(n1140), .Y(n1143) );
  INVX2TS U716 ( .A(n686), .Y(n1205) );
  CLKAND2X2TS U717 ( .A(n1255), .B(n1254), .Y(n1249) );
  MXI2XLTS U718 ( .A(n1146), .B(n1145), .S0(n1286), .Y(n1207) );
  MXI2XLTS U719 ( .A(n1173), .B(n1172), .S0(n1292), .Y(n1206) );
  MXI2XLTS U720 ( .A(n1215), .B(n1214), .S0(n1266), .Y(n1239) );
  MXI2XLTS U721 ( .A(n1210), .B(n1209), .S0(n1196), .Y(n1242) );
  INVX2TS U722 ( .A(n1208), .Y(n1209) );
  MXI2XLTS U723 ( .A(n1212), .B(n1211), .S0(n1225), .Y(n1241) );
  INVX2TS U724 ( .A(n1243), .Y(n1247) );
  INVX2TS U725 ( .A(n1256), .Y(n690) );
  INVX2TS U726 ( .A(n704), .Y(n692) );
  XOR2XLTS U727 ( .A(sumIn[47]), .B(n707), .Y(n777) );
  INVX2TS U728 ( .A(n902), .Y(n843) );
  INVX2TS U729 ( .A(n1283), .Y(n1101) );
  INVX2TS U730 ( .A(n1173), .Y(n1119) );
  MXI2XLTS U731 ( .A(n1053), .B(n1083), .S0(n1091), .Y(n1142) );
  MXI2XLTS U732 ( .A(n1085), .B(n1084), .S0(n1095), .Y(n1140) );
  MXI2XLTS U733 ( .A(n1087), .B(n1086), .S0(n1091), .Y(n1172) );
  AO21XLTS U734 ( .A0(n1172), .A1(n1119), .B0(n1116), .Y(n1117) );
  MXI2XLTS U735 ( .A(n1080), .B(n1079), .S0(n1101), .Y(n1135) );
  INVX2TS U736 ( .A(n1078), .Y(n1079) );
  MXI2XLTS U737 ( .A(n1082), .B(n1081), .S0(n1108), .Y(n1136) );
  INVX2TS U738 ( .A(n1284), .Y(n1108) );
  XOR2XLTS U739 ( .A(sumIn[87]), .B(n993), .Y(n1070) );
  INVX2TS U740 ( .A(n1082), .Y(n1058) );
  XOR2XLTS U741 ( .A(n1062), .B(sumIn[98]), .Y(n1076) );
  XOR2XLTS U742 ( .A(sumIn[67]), .B(n916), .Y(n990) );
  INVX2TS U743 ( .A(n1138), .Y(n899) );
  INVX2TS U744 ( .A(n1147), .Y(n892) );
  MXI2XLTS U745 ( .A(n797), .B(n868), .S0(n1287), .Y(n1145) );
  NAND2BXLTS U746 ( .AN(n894), .B(n1146), .Y(n897) );
  MXI2XLTS U747 ( .A(n866), .B(n865), .S0(n1288), .Y(n1139) );
  MXI2XLTS U748 ( .A(n861), .B(n860), .S0(n859), .Y(n1182) );
  INVX2TS U749 ( .A(n858), .Y(n861) );
  MXI2XLTS U750 ( .A(n902), .B(n901), .S0(n900), .Y(n1181) );
  XOR2XLTS U751 ( .A(sumIn[27]), .B(n780), .Y(n852) );
  XOR2XLTS U752 ( .A(n787), .B(sumIn[38]), .Y(n856) );
  INVX2TS U753 ( .A(n1197), .Y(n1189) );
  OAI31X1TS U754 ( .A0(n1187), .A1(n1201), .A2(n1185), .B0(n1184), .Y(n1186)
         );
  INVX2TS U755 ( .A(n1183), .Y(n1185) );
  NOR3BXLTS U756 ( .AN(n711), .B(sumIn[48]), .C(n722), .Y(n715) );
  NOR3BXLTS U757 ( .AN(n713), .B(sumIn[58]), .C(n730), .Y(n773) );
  NOR3BXLTS U758 ( .AN(n784), .B(sumIn[28]), .C(n795), .Y(n788) );
  NOR3BXLTS U759 ( .AN(n786), .B(sumIn[38]), .C(n803), .Y(n848) );
  NOR3BXLTS U760 ( .AN(n987), .B(sumIn[78]), .C(n921), .Y(n1071) );
  NAND3BXLTS U761 ( .AN(sumIn[68]), .B(n986), .C(n985), .Y(n1072) );
  NOR3BXLTS U762 ( .AN(n1067), .B(sumIn[98]), .C(n998), .Y(n1126) );
  NAND3BXLTS U763 ( .AN(sumIn[88]), .B(n1066), .C(n1065), .Y(n1125) );
  MXI2XLTS U764 ( .A(n777), .B(n776), .S0(n859), .Y(n913) );
  INVX2TS U765 ( .A(n771), .Y(n776) );
  MXI2XLTS U766 ( .A(n990), .B(n989), .S0(n1101), .Y(n1130) );
  INVX2TS U767 ( .A(n981), .Y(n989) );
  MXI2XLTS U768 ( .A(n1204), .B(n1203), .S0(n1266), .Y(n1255) );
  INVX2TS U769 ( .A(n1202), .Y(n1203) );
  MXI2XLTS U770 ( .A(n1205), .B(n685), .S0(n1225), .Y(n1254) );
  OAI31X1TS U771 ( .A0(n1251), .A1(n1252), .A2(n1249), .B0(n1248), .Y(n1250)
         );
  MXI2XLTS U772 ( .A(n1207), .B(n1206), .S0(n1196), .Y(n1252) );
  OAI31X1TS U773 ( .A0(n639), .A1(n638), .A2(n656), .B0(n637), .Y(n1257) );
  XOR2XLTS U774 ( .A(n635), .B(sumIn[6]), .Y(n1256) );
  MXI2XLTS U775 ( .A(n1137), .B(n1136), .S0(n1141), .Y(n1201) );
  INVX2TS U776 ( .A(n1135), .Y(n1137) );
  MXI2XLTS U777 ( .A(n1182), .B(n1181), .S0(n1180), .Y(n1200) );
  INVX2TS U778 ( .A(n856), .Y(n847) );
  MXI2XLTS U779 ( .A(n1075), .B(n1074), .S0(n1101), .Y(n1131) );
  INVX2TS U780 ( .A(n1073), .Y(n1075) );
  MXI2XLTS U781 ( .A(n1077), .B(n1076), .S0(n1108), .Y(n1132) );
  INVX2TS U782 ( .A(n1130), .Y(n1123) );
  MXI2XLTS U783 ( .A(n1070), .B(n1069), .S0(n1108), .Y(n1129) );
  INVX2TS U784 ( .A(n1060), .Y(n1069) );
  AO21XLTS U785 ( .A0(n1068), .A1(n1125), .B0(n1126), .Y(n602) );
  INVX2TS U786 ( .A(n1076), .Y(n1063) );
  AO21XLTS U787 ( .A0(n988), .A1(n1072), .B0(n1071), .Y(n601) );
  INVX2TS U788 ( .A(n1182), .Y(n904) );
  MXI2XLTS U789 ( .A(n852), .B(n851), .S0(n862), .Y(n912) );
  INVX2TS U790 ( .A(n845), .Y(n851) );
  INVX2TS U791 ( .A(n913), .Y(n905) );
  MXI2XLTS U792 ( .A(n857), .B(n856), .S0(n862), .Y(n1133) );
  MXI2XLTS U793 ( .A(n855), .B(n854), .S0(n859), .Y(n1134) );
  INVX2TS U794 ( .A(n853), .Y(n855) );
  INVX2TS U795 ( .A(n1281), .Y(n1194) );
  NAND2BXLTS U796 ( .AN(n1126), .B(n1125), .Y(n1192) );
  NAND2BXLTS U797 ( .AN(n1134), .B(n1133), .Y(n1268) );
  OAI31X1TS U798 ( .A0(n694), .A1(n693), .A2(n695), .B0(n628), .Y(n703) );
  OAI31X1TS U799 ( .A0(n630), .A1(n629), .A2(n633), .B0(n620), .Y(n704) );
  MXI2XLTS U800 ( .A(n913), .B(n912), .S0(n1164), .Y(n1198) );
  MXI2XLTS U801 ( .A(n1130), .B(n1129), .S0(n1141), .Y(n1197) );
  MX2X1TS U802 ( .A(n1201), .B(n1200), .S0(n1195), .Y(n1260) );
  MXI2XLTS U803 ( .A(n1257), .B(n1256), .S0(n702), .Y(n1258) );
  NAND2BXLTS U804 ( .AN(n1192), .B(n1191), .Y(n1279) );
  NOR3BXLTS U805 ( .AN(n700), .B(sumIn[18]), .C(n699), .Y(n1276) );
  NAND3BXLTS U806 ( .AN(sumIn[8]), .B(n698), .C(n631), .Y(n1275) );
  MXI2XLTS U807 ( .A(n1268), .B(n1267), .S0(n1266), .Y(n1273) );
  INVX2TS U808 ( .A(n1265), .Y(n1267) );
  OAI21XLTS U809 ( .A0(n1264), .A1(n1263), .B0(n1262), .Y(n1274) );
  MXI2XLTS U810 ( .A(n1198), .B(n1197), .S0(n1199), .Y(n1263) );
  MXI2XLTS U811 ( .A(n704), .B(n703), .S0(n1225), .Y(n1264) );
  INVX2TS U812 ( .A(n1277), .Y(n1278) );
  NAND2BXLTS U813 ( .AN(n1276), .B(n1275), .Y(n1277) );
  OAI31X1TS U814 ( .A0(n1013), .A1(n1012), .A2(n1023), .B0(n1011), .Y(n1019)
         );
  INVX2TS U815 ( .A(n1019), .Y(n1053) );
  OAI31X1TS U816 ( .A0(n936), .A1(n935), .A2(n945), .B0(n934), .Y(n1085) );
  INVX2TS U817 ( .A(n1085), .Y(n976) );
  OAI31X1TS U818 ( .A0(n727), .A1(n726), .A2(n730), .B0(n725), .Y(n865) );
  INVX2TS U819 ( .A(n865), .Y(n766) );
  OAI31X1TS U820 ( .A0(n800), .A1(n799), .A2(n803), .B0(n798), .Y(n863) );
  INVX2TS U821 ( .A(n863), .Y(n839) );
  INVX2TS U822 ( .A(n1294), .Y(n1196) );
  OAI31X1TS U823 ( .A0(n644), .A1(n643), .A2(n699), .B0(n642), .Y(n651) );
  INVX2TS U824 ( .A(n651), .Y(n685) );
  AOI21X1TS U825 ( .A0(n850), .A1(n849), .B0(n848), .Y(n599) );
  AOI21X1TS U826 ( .A0(n775), .A1(n774), .B0(n773), .Y(n600) );
  INVX2TS U827 ( .A(n985), .Y(n924) );
  INVX2TS U828 ( .A(n1065), .Y(n1001) );
  INVX2TS U829 ( .A(sumIn[53]), .Y(n603) );
  INVX2TS U830 ( .A(n603), .Y(n739) );
  INVX2TS U831 ( .A(sumIn[52]), .Y(n604) );
  INVX2TS U832 ( .A(n604), .Y(n745) );
  INVX2TS U833 ( .A(sumIn[51]), .Y(n736) );
  INVX2TS U834 ( .A(n736), .Y(n754) );
  INVX2TS U835 ( .A(sumIn[50]), .Y(n752) );
  INVX2TS U836 ( .A(n752), .Y(n751) );
  NOR4XLTS U837 ( .A(n739), .B(n745), .C(n754), .D(n751), .Y(n733) );
  INVX2TS U838 ( .A(sumIn[54]), .Y(n605) );
  INVX2TS U839 ( .A(n605), .Y(n732) );
  NOR2BX1TS U840 ( .AN(n733), .B(n732), .Y(n727) );
  INVX2TS U841 ( .A(sumIn[55]), .Y(n606) );
  INVX2TS U842 ( .A(n606), .Y(n726) );
  NOR2BX1TS U843 ( .AN(n727), .B(n726), .Y(n720) );
  NOR2XLTS U844 ( .A(sumIn[57]), .B(n708), .Y(n713) );
  INVX2TS U845 ( .A(sumIn[59]), .Y(n607) );
  INVX2TS U846 ( .A(n607), .Y(n753) );
  CLKBUFX2TS U847 ( .A(n753), .Y(n718) );
  INVX2TS U848 ( .A(n718), .Y(n730) );
  INVX2TS U849 ( .A(sumIn[42]), .Y(n608) );
  INVX2TS U850 ( .A(n608), .Y(n744) );
  INVX2TS U851 ( .A(sumIn[41]), .Y(n609) );
  INVX2TS U852 ( .A(n609), .Y(n750) );
  INVX2TS U853 ( .A(sumIn[40]), .Y(n748) );
  INVX2TS U854 ( .A(n748), .Y(n742) );
  NOR4XLTS U855 ( .A(sumIn[43]), .B(n744), .C(n750), .D(n742), .Y(n723) );
  NOR2XLTS U856 ( .A(sumIn[45]), .B(n728), .Y(n716) );
  NOR2XLTS U857 ( .A(sumIn[47]), .B(n706), .Y(n711) );
  INVX2TS U858 ( .A(sumIn[49]), .Y(n705) );
  INVX2TS U859 ( .A(n705), .Y(n741) );
  CLKBUFX2TS U860 ( .A(n741), .Y(n710) );
  NOR2XLTS U861 ( .A(n773), .B(n715), .Y(n909) );
  INVX2TS U862 ( .A(sumIn[33]), .Y(n610) );
  INVX2TS U863 ( .A(n610), .Y(n812) );
  INVX2TS U864 ( .A(sumIn[32]), .Y(n611) );
  INVX2TS U865 ( .A(n611), .Y(n818) );
  INVX2TS U866 ( .A(sumIn[31]), .Y(n809) );
  INVX2TS U867 ( .A(n809), .Y(n827) );
  INVX2TS U868 ( .A(sumIn[30]), .Y(n825) );
  INVX2TS U869 ( .A(n825), .Y(n822) );
  NOR4XLTS U870 ( .A(n812), .B(n818), .C(n827), .D(n822), .Y(n806) );
  INVX2TS U871 ( .A(sumIn[34]), .Y(n612) );
  INVX2TS U872 ( .A(n612), .Y(n805) );
  NOR2BX1TS U873 ( .AN(n806), .B(n805), .Y(n800) );
  INVX2TS U874 ( .A(sumIn[35]), .Y(n613) );
  INVX2TS U875 ( .A(n613), .Y(n799) );
  NOR2BX1TS U876 ( .AN(n800), .B(n799), .Y(n793) );
  NOR2XLTS U877 ( .A(sumIn[37]), .B(n781), .Y(n786) );
  INVX2TS U878 ( .A(sumIn[39]), .Y(n614) );
  INVX2TS U879 ( .A(n614), .Y(n826) );
  CLKBUFX2TS U880 ( .A(n826), .Y(n791) );
  INVX2TS U881 ( .A(n791), .Y(n803) );
  INVX2TS U882 ( .A(sumIn[21]), .Y(n615) );
  INVX2TS U883 ( .A(n615), .Y(n824) );
  INVX2TS U884 ( .A(sumIn[20]), .Y(n821) );
  INVX2TS U885 ( .A(n821), .Y(n815) );
  INVX2TS U886 ( .A(sumIn[22]), .Y(n616) );
  INVX2TS U887 ( .A(n616), .Y(n817) );
  NOR4XLTS U888 ( .A(n824), .B(n815), .C(sumIn[23]), .D(n817), .Y(n796) );
  NOR2XLTS U889 ( .A(sumIn[25]), .B(n801), .Y(n789) );
  NOR2XLTS U890 ( .A(sumIn[27]), .B(n779), .Y(n784) );
  INVX2TS U891 ( .A(sumIn[29]), .Y(n778) );
  INVX2TS U892 ( .A(n778), .Y(n814) );
  CLKBUFX2TS U893 ( .A(n814), .Y(n783) );
  NOR2XLTS U894 ( .A(n848), .B(n788), .Y(n908) );
  NAND2X1TS U895 ( .A(n909), .B(n908), .Y(n1281) );
  INVX2TS U896 ( .A(sumIn[2]), .Y(n617) );
  INVX2TS U897 ( .A(n617), .Y(n662) );
  INVX2TS U898 ( .A(sumIn[1]), .Y(n618) );
  INVX2TS U899 ( .A(n618), .Y(n668) );
  INVX2TS U900 ( .A(sumIn[0]), .Y(n666) );
  INVX2TS U901 ( .A(n666), .Y(n660) );
  NOR4XLTS U902 ( .A(sumIn[3]), .B(n662), .C(n668), .D(n660), .Y(n641) );
  NOR2XLTS U903 ( .A(sumIn[5]), .B(n646), .Y(n634) );
  NOR2BX1TS U904 ( .AN(n634), .B(sumIn[6]), .Y(n630) );
  INVX2TS U905 ( .A(sumIn[7]), .Y(n619) );
  INVX2TS U906 ( .A(n619), .Y(n629) );
  INVX2TS U907 ( .A(sumIn[9]), .Y(n645) );
  INVX2TS U908 ( .A(n645), .Y(n659) );
  CLKBUFX2TS U909 ( .A(n659), .Y(n631) );
  INVX2TS U910 ( .A(n631), .Y(n633) );
  OAI21XLTS U911 ( .A0(n630), .A1(n633), .B0(n629), .Y(n620) );
  INVX2TS U912 ( .A(sumIn[13]), .Y(n621) );
  INVX2TS U913 ( .A(n621), .Y(n657) );
  INVX2TS U914 ( .A(sumIn[12]), .Y(n622) );
  INVX2TS U915 ( .A(n622), .Y(n663) );
  INVX2TS U916 ( .A(sumIn[11]), .Y(n654) );
  INVX2TS U917 ( .A(n654), .Y(n672) );
  INVX2TS U918 ( .A(sumIn[10]), .Y(n670) );
  INVX2TS U919 ( .A(n670), .Y(n669) );
  NOR4XLTS U920 ( .A(n657), .B(n663), .C(n672), .D(n669), .Y(n650) );
  INVX2TS U921 ( .A(sumIn[14]), .Y(n623) );
  INVX2TS U922 ( .A(n623), .Y(n649) );
  NOR2BX1TS U923 ( .AN(n650), .B(n649), .Y(n644) );
  INVX2TS U924 ( .A(sumIn[15]), .Y(n624) );
  INVX2TS U925 ( .A(n624), .Y(n643) );
  NOR2BX1TS U926 ( .AN(n644), .B(n643), .Y(n639) );
  INVX2TS U927 ( .A(sumIn[16]), .Y(n625) );
  INVX2TS U928 ( .A(n625), .Y(n638) );
  NOR2BX1TS U929 ( .AN(n639), .B(n638), .Y(n694) );
  INVX2TS U930 ( .A(sumIn[17]), .Y(n626) );
  INVX2TS U931 ( .A(n626), .Y(n693) );
  INVX2TS U932 ( .A(sumIn[19]), .Y(n627) );
  INVX2TS U933 ( .A(n627), .Y(n671) );
  CLKBUFX2TS U934 ( .A(n671), .Y(n636) );
  INVX2TS U935 ( .A(n636), .Y(n695) );
  INVX2TS U936 ( .A(n636), .Y(n656) );
  OAI21XLTS U937 ( .A0(n694), .A1(n656), .B0(n693), .Y(n628) );
  NOR2BX1TS U938 ( .AN(n630), .B(n629), .Y(n698) );
  OAI21XLTS U939 ( .A0(n698), .A1(n633), .B0(sumIn[8]), .Y(n632) );
  OAI21XLTS U940 ( .A0(sumIn[8]), .A1(n633), .B0(n632), .Y(n1269) );
  NOR2XLTS U941 ( .A(n645), .B(n634), .Y(n635) );
  INVX2TS U942 ( .A(n636), .Y(n699) );
  OAI21XLTS U943 ( .A0(n639), .A1(n699), .B0(n638), .Y(n637) );
  OAI21XLTS U944 ( .A0(n641), .A1(n645), .B0(sumIn[4]), .Y(n640) );
  OAI31XLTS U945 ( .A0(n641), .A1(sumIn[4]), .A2(n645), .B0(n640), .Y(n1243)
         );
  OAI21XLTS U946 ( .A0(n644), .A1(n695), .B0(n643), .Y(n642) );
  NAND2X1TS U947 ( .A(n646), .B(n659), .Y(n647) );
  XNOR2X1TS U948 ( .A(sumIn[5]), .B(n647), .Y(n686) );
  OAI21XLTS U949 ( .A0(n650), .A1(n656), .B0(n649), .Y(n648) );
  AOI21X1TS U950 ( .A0(n651), .A1(n1205), .B0(n1244), .Y(n652) );
  NAND2X1TS U951 ( .A(n1243), .B(n652), .Y(n688) );
  NAND2X1TS U952 ( .A(n1243), .B(n686), .Y(n683) );
  AOI21X1TS U953 ( .A0(n1243), .A1(n685), .B0(n652), .Y(n682) );
  XNOR2X1TS U954 ( .A(sumIn[3]), .B(n653), .Y(n1212) );
  INVX2TS U955 ( .A(n654), .Y(n674) );
  NOR3XLTS U956 ( .A(n663), .B(n674), .C(n669), .Y(n658) );
  OAI21XLTS U957 ( .A0(n658), .A1(n699), .B0(n657), .Y(n655) );
  OAI21XLTS U958 ( .A0(n668), .A1(n660), .B0(n659), .Y(n661) );
  XNOR2X1TS U959 ( .A(n662), .B(n661), .Y(n1231) );
  OAI21XLTS U960 ( .A0(n674), .A1(n669), .B0(n671), .Y(n664) );
  OAI2BB2XLTS U961 ( .B0(n1211), .B1(n677), .A0N(n1231), .A1N(n1234), .Y(n665)
         );
  OAI2BB1X1TS U962 ( .A0N(n677), .A1N(n1211), .B0(n665), .Y(n681) );
  INVX2TS U963 ( .A(n666), .Y(n1216) );
  NAND2X1TS U964 ( .A(n631), .B(n1216), .Y(n667) );
  XNOR2X1TS U965 ( .A(n668), .B(n667), .Y(n1227) );
  INVX2TS U966 ( .A(n670), .Y(n1217) );
  NAND2X1TS U967 ( .A(n671), .B(n1217), .Y(n673) );
  XNOR2X1TS U968 ( .A(n673), .B(n672), .Y(n1226) );
  AOI222XLTS U969 ( .A0(n676), .A1(n675), .B0(n676), .B1(n674), .C0(n675), 
        .C1(n1226), .Y(n679) );
  NAND2X1TS U970 ( .A(n1211), .B(n677), .Y(n678) );
  OAI211XLTS U971 ( .A0(n1231), .A1(n1234), .B0(n679), .C0(n678), .Y(n680) );
  AOI22X1TS U972 ( .A0(n683), .A1(n682), .B0(n681), .B1(n680), .Y(n684) );
  AOI21X1TS U973 ( .A0(n686), .A1(n685), .B0(n684), .Y(n687) );
  OAI211XLTS U974 ( .A0(n1257), .A1(n690), .B0(n688), .C0(n687), .Y(n689) );
  OAI2BB1X1TS U975 ( .A0N(n690), .A1N(n1257), .B0(n689), .Y(n691) );
  AOI222XLTS U976 ( .A0(n703), .A1(n692), .B0(n703), .B1(n691), .C0(n692), 
        .C1(n691), .Y(n697) );
  NOR2BX1TS U977 ( .AN(n694), .B(n693), .Y(n700) );
  NOR2XLTS U978 ( .A(n695), .B(n700), .Y(n696) );
  XNOR2X1TS U979 ( .A(n696), .B(sumIn[18]), .Y(n1270) );
  AOI222XLTS U980 ( .A0(n1269), .A1(n697), .B0(n1269), .B1(n1270), .C0(n697), 
        .C1(n1270), .Y(n701) );
  AOI21X1TS U981 ( .A0(n701), .A1(n1275), .B0(n1276), .Y(n702) );
  INVX2TS U982 ( .A(n702), .Y(n1225) );
  NAND2X1TS U983 ( .A(n706), .B(n710), .Y(n707) );
  NAND2X1TS U984 ( .A(n708), .B(n753), .Y(n709) );
  XNOR2X1TS U985 ( .A(sumIn[57]), .B(n709), .Y(n771) );
  INVX2TS U986 ( .A(n710), .Y(n722) );
  OAI21XLTS U987 ( .A0(n711), .A1(n705), .B0(sumIn[48]), .Y(n712) );
  OAI21XLTS U988 ( .A0(sumIn[48]), .A1(n722), .B0(n712), .Y(n853) );
  NOR2XLTS U989 ( .A(n730), .B(n713), .Y(n714) );
  XNOR2X1TS U990 ( .A(n714), .B(sumIn[58]), .Y(n854) );
  AOI21X1TS U991 ( .A0(n853), .A1(n854), .B0(n715), .Y(n775) );
  NOR2XLTS U992 ( .A(n722), .B(n716), .Y(n717) );
  XNOR2X1TS U993 ( .A(n717), .B(sumIn[46]), .Y(n858) );
  INVX2TS U994 ( .A(n718), .Y(n737) );
  OAI21XLTS U995 ( .A0(n720), .A1(n737), .B0(sumIn[56]), .Y(n719) );
  OAI31XLTS U996 ( .A0(n720), .A1(sumIn[56]), .A2(n607), .B0(n719), .Y(n860)
         );
  OAI21XLTS U997 ( .A0(n723), .A1(n705), .B0(sumIn[44]), .Y(n721) );
  OAI31XLTS U998 ( .A0(n723), .A1(sumIn[44]), .A2(n722), .B0(n721), .Y(n724)
         );
  OAI21XLTS U999 ( .A0(n727), .A1(n607), .B0(n726), .Y(n725) );
  NAND2X1TS U1000 ( .A(n728), .B(n741), .Y(n729) );
  XNOR2X1TS U1001 ( .A(sumIn[45]), .B(n729), .Y(n866) );
  OAI21XLTS U1002 ( .A0(n733), .A1(n730), .B0(n732), .Y(n731) );
  NAND2X1TS U1003 ( .A(n724), .B(n734), .Y(n768) );
  NAND2X1TS U1004 ( .A(n724), .B(n866), .Y(n764) );
  AOI21X1TS U1005 ( .A0(n724), .A1(n766), .B0(n734), .Y(n763) );
  INVX2TS U1006 ( .A(n736), .Y(n756) );
  NOR3XLTS U1007 ( .A(n745), .B(n756), .C(n751), .Y(n740) );
  OAI21XLTS U1008 ( .A0(n740), .A1(n737), .B0(n739), .Y(n738) );
  OAI21XLTS U1009 ( .A0(n750), .A1(n742), .B0(n741), .Y(n743) );
  XNOR2X1TS U1010 ( .A(n744), .B(n743), .Y(n877) );
  OAI21XLTS U1011 ( .A0(n756), .A1(n751), .B0(n753), .Y(n746) );
  OAI2BB2XLTS U1012 ( .B0(n869), .B1(n871), .A0N(n877), .A1N(n875), .Y(n747)
         );
  OAI2BB1X1TS U1013 ( .A0N(n871), .A1N(n869), .B0(n747), .Y(n762) );
  INVX2TS U1014 ( .A(n748), .Y(n886) );
  NAND2X1TS U1015 ( .A(n710), .B(n886), .Y(n749) );
  XNOR2X1TS U1016 ( .A(n750), .B(n749), .Y(n881) );
  INVX2TS U1017 ( .A(n752), .Y(n885) );
  NAND2X1TS U1018 ( .A(n753), .B(n885), .Y(n755) );
  XNOR2X1TS U1019 ( .A(n755), .B(n754), .Y(n880) );
  AOI222XLTS U1020 ( .A0(n758), .A1(n757), .B0(n758), .B1(n756), .C0(n757), 
        .C1(n880), .Y(n760) );
  NAND2X1TS U1021 ( .A(n869), .B(n871), .Y(n759) );
  OAI211XLTS U1022 ( .A0(n877), .A1(n875), .B0(n760), .C0(n759), .Y(n761) );
  AOI22X1TS U1023 ( .A0(n764), .A1(n763), .B0(n762), .B1(n761), .Y(n765) );
  AOI21X1TS U1024 ( .A0(n866), .A1(n766), .B0(n765), .Y(n767) );
  OAI211XLTS U1025 ( .A0(n860), .A1(n858), .B0(n768), .C0(n767), .Y(n769) );
  OAI2BB1X1TS U1026 ( .A0N(n858), .A1N(n860), .B0(n769), .Y(n770) );
  AOI222XLTS U1027 ( .A0(n771), .A1(n777), .B0(n771), .B1(n770), .C0(n777), 
        .C1(n770), .Y(n772) );
  OAI21XLTS U1028 ( .A0(n853), .A1(n854), .B0(n772), .Y(n774) );
  INVX2TS U1029 ( .A(n600), .Y(n859) );
  NAND2X1TS U1030 ( .A(n779), .B(n783), .Y(n780) );
  NAND2X1TS U1031 ( .A(n781), .B(n826), .Y(n782) );
  XNOR2X1TS U1032 ( .A(sumIn[37]), .B(n782), .Y(n845) );
  INVX2TS U1033 ( .A(n783), .Y(n795) );
  OAI21XLTS U1034 ( .A0(n784), .A1(n778), .B0(sumIn[28]), .Y(n785) );
  OAI21XLTS U1035 ( .A0(sumIn[28]), .A1(n795), .B0(n785), .Y(n857) );
  NOR2XLTS U1036 ( .A(n803), .B(n786), .Y(n787) );
  AOI21X1TS U1037 ( .A0(n857), .A1(n847), .B0(n788), .Y(n850) );
  NOR2XLTS U1038 ( .A(n795), .B(n789), .Y(n790) );
  INVX2TS U1039 ( .A(n791), .Y(n810) );
  OAI21XLTS U1040 ( .A0(n793), .A1(n810), .B0(sumIn[36]), .Y(n792) );
  OAI31XLTS U1041 ( .A0(n793), .A1(sumIn[36]), .A2(n614), .B0(n792), .Y(n901)
         );
  OAI21XLTS U1042 ( .A0(n796), .A1(n778), .B0(sumIn[24]), .Y(n794) );
  OAI31XLTS U1043 ( .A0(n796), .A1(sumIn[24]), .A2(n795), .B0(n794), .Y(n797)
         );
  OAI21XLTS U1044 ( .A0(n800), .A1(n614), .B0(n799), .Y(n798) );
  NAND2X1TS U1045 ( .A(n801), .B(n814), .Y(n802) );
  XNOR2X1TS U1046 ( .A(sumIn[25]), .B(n802), .Y(n864) );
  OAI21XLTS U1047 ( .A0(n806), .A1(n803), .B0(n805), .Y(n804) );
  NAND2X1TS U1048 ( .A(n797), .B(n807), .Y(n841) );
  NAND2X1TS U1049 ( .A(n797), .B(n864), .Y(n837) );
  AOI21X1TS U1050 ( .A0(n797), .A1(n839), .B0(n807), .Y(n836) );
  INVX2TS U1051 ( .A(n809), .Y(n829) );
  NOR3XLTS U1052 ( .A(n818), .B(n829), .C(n822), .Y(n813) );
  OAI21XLTS U1053 ( .A0(n813), .A1(n810), .B0(n812), .Y(n811) );
  OAI21XLTS U1054 ( .A0(n824), .A1(n815), .B0(n814), .Y(n816) );
  XNOR2X1TS U1055 ( .A(n817), .B(n816), .Y(n872) );
  OAI21XLTS U1056 ( .A0(n829), .A1(n822), .B0(n826), .Y(n819) );
  OAI2BB2XLTS U1057 ( .B0(n889), .B1(n891), .A0N(n872), .A1N(n873), .Y(n820)
         );
  OAI2BB1X1TS U1058 ( .A0N(n891), .A1N(n889), .B0(n820), .Y(n835) );
  INVX2TS U1059 ( .A(n821), .Y(n879) );
  NAND2X1TS U1060 ( .A(n783), .B(n879), .Y(n823) );
  INVX2TS U1061 ( .A(n825), .Y(n878) );
  NAND2X1TS U1062 ( .A(n826), .B(n878), .Y(n828) );
  AOI222XLTS U1063 ( .A0(n831), .A1(n883), .B0(n831), .B1(n830), .C0(n883), 
        .C1(n829), .Y(n833) );
  NAND2X1TS U1064 ( .A(n889), .B(n891), .Y(n832) );
  OAI211XLTS U1065 ( .A0(n872), .A1(n873), .B0(n833), .C0(n832), .Y(n834) );
  AOI22X1TS U1066 ( .A0(n837), .A1(n836), .B0(n835), .B1(n834), .Y(n838) );
  AOI21X1TS U1067 ( .A0(n864), .A1(n839), .B0(n838), .Y(n840) );
  OAI211XLTS U1068 ( .A0(n901), .A1(n843), .B0(n841), .C0(n840), .Y(n842) );
  OAI2BB1X1TS U1069 ( .A0N(n843), .A1N(n901), .B0(n842), .Y(n844) );
  AOI222XLTS U1070 ( .A0(n845), .A1(n852), .B0(n845), .B1(n844), .C0(n852), 
        .C1(n844), .Y(n846) );
  OAI21XLTS U1071 ( .A0(n857), .A1(n847), .B0(n846), .Y(n849) );
  INVX2TS U1072 ( .A(n599), .Y(n862) );
  INVX2TS U1073 ( .A(n600), .Y(n1288) );
  NOR2XLTS U1074 ( .A(n1139), .B(n899), .Y(n894) );
  INVX2TS U1075 ( .A(n600), .Y(n884) );
  INVX2TS U1076 ( .A(n599), .Y(n1287) );
  INVX2TS U1077 ( .A(n599), .Y(n900) );
  OAI21XLTS U1078 ( .A0(n1156), .A1(n1154), .B0(n1161), .Y(n887) );
  OAI2BB2XLTS U1079 ( .B0(n1160), .B1(n887), .A0N(n1156), .A1N(n1154), .Y(n888) );
  AOI222XLTS U1080 ( .A0(n1163), .A1(n1166), .B0(n1163), .B1(n888), .C0(n1166), 
        .C1(n888), .Y(n893) );
  AOI222XLTS U1081 ( .A0(n1148), .A1(n893), .B0(n1148), .B1(n892), .C0(n893), 
        .C1(n892), .Y(n896) );
  OAI21XLTS U1082 ( .A0(n1145), .A1(n894), .B0(n897), .Y(n895) );
  OAI2BB2XLTS U1083 ( .B0(n897), .B1(n1145), .A0N(n896), .A1N(n895), .Y(n898)
         );
  AOI21X1TS U1084 ( .A0(n899), .A1(n1139), .B0(n898), .Y(n903) );
  AOI222XLTS U1085 ( .A0(n904), .A1(n903), .B0(n904), .B1(n1181), .C0(n903), 
        .C1(n1181), .Y(n906) );
  AOI222XLTS U1086 ( .A0(n912), .A1(n906), .B0(n912), .B1(n905), .C0(n906), 
        .C1(n905), .Y(n907) );
  AOI21X1TS U1087 ( .A0(n1134), .A1(n1133), .B0(n907), .Y(n911) );
  OAI21XLTS U1088 ( .A0(n1134), .A1(n1133), .B0(n908), .Y(n910) );
  OAI21XLTS U1089 ( .A0(n911), .A1(n910), .B0(n909), .Y(n1293) );
  CLKBUFX2TS U1090 ( .A(n1293), .Y(n1144) );
  INVX2TS U1091 ( .A(n1144), .Y(n1164) );
  INVX2TS U1092 ( .A(sumIn[61]), .Y(n914) );
  INVX2TS U1093 ( .A(n914), .Y(n960) );
  INVX2TS U1094 ( .A(sumIn[60]), .Y(n956) );
  INVX2TS U1095 ( .A(n956), .Y(n950) );
  INVX2TS U1096 ( .A(sumIn[62]), .Y(n915) );
  INVX2TS U1097 ( .A(n915), .Y(n952) );
  NOR4XLTS U1098 ( .A(n960), .B(n950), .C(sumIn[63]), .D(n952), .Y(n932) );
  NOR2XLTS U1099 ( .A(sumIn[65]), .B(n937), .Y(n927) );
  INVX2TS U1100 ( .A(sumIn[69]), .Y(n923) );
  INVX2TS U1101 ( .A(n923), .Y(n958) );
  NAND2X1TS U1102 ( .A(n925), .B(n958), .Y(n916) );
  INVX2TS U1103 ( .A(sumIn[73]), .Y(n917) );
  INVX2TS U1104 ( .A(n917), .Y(n948) );
  INVX2TS U1105 ( .A(sumIn[72]), .Y(n918) );
  INVX2TS U1106 ( .A(n918), .Y(n953) );
  INVX2TS U1107 ( .A(sumIn[71]), .Y(n944) );
  INVX2TS U1108 ( .A(n944), .Y(n963) );
  INVX2TS U1109 ( .A(sumIn[70]), .Y(n961) );
  INVX2TS U1110 ( .A(n961), .Y(n957) );
  NOR4XLTS U1111 ( .A(n948), .B(n953), .C(n963), .D(n957), .Y(n941) );
  INVX2TS U1112 ( .A(sumIn[74]), .Y(n919) );
  INVX2TS U1113 ( .A(n919), .Y(n940) );
  NOR2BX1TS U1114 ( .AN(n941), .B(n940), .Y(n936) );
  INVX2TS U1115 ( .A(sumIn[75]), .Y(n920) );
  INVX2TS U1116 ( .A(n920), .Y(n935) );
  NOR2BX1TS U1117 ( .AN(n936), .B(n935), .Y(n930) );
  INVX2TS U1118 ( .A(sumIn[79]), .Y(n921) );
  INVX2TS U1119 ( .A(n921), .Y(n962) );
  NAND2X1TS U1120 ( .A(n982), .B(n962), .Y(n922) );
  XNOR2X1TS U1121 ( .A(sumIn[77]), .B(n922), .Y(n981) );
  INVX2TS U1122 ( .A(n923), .Y(n985) );
  NOR2XLTS U1123 ( .A(sumIn[67]), .B(n925), .Y(n986) );
  OAI21XLTS U1124 ( .A0(n986), .A1(n924), .B0(sumIn[68]), .Y(n926) );
  OAI21XLTS U1125 ( .A0(sumIn[68]), .A1(n924), .B0(n926), .Y(n1073) );
  NOR2XLTS U1126 ( .A(n923), .B(n927), .Y(n928) );
  XNOR2X1TS U1127 ( .A(n928), .B(sumIn[66]), .Y(n1080) );
  CLKBUFX2TS U1128 ( .A(n962), .Y(n933) );
  INVX2TS U1129 ( .A(n933), .Y(n947) );
  INVX2TS U1130 ( .A(n933), .Y(n945) );
  OAI21XLTS U1131 ( .A0(n930), .A1(n945), .B0(sumIn[76]), .Y(n929) );
  OAI31XLTS U1132 ( .A0(n930), .A1(sumIn[76]), .A2(n947), .B0(n929), .Y(n1078)
         );
  OAI21XLTS U1133 ( .A0(n932), .A1(n924), .B0(sumIn[64]), .Y(n931) );
  OAI31XLTS U1134 ( .A0(n932), .A1(sumIn[64]), .A2(n924), .B0(n931), .Y(n1088)
         );
  OAI21XLTS U1135 ( .A0(n936), .A1(n947), .B0(n935), .Y(n934) );
  NAND2X1TS U1136 ( .A(n937), .B(n958), .Y(n938) );
  XNOR2X1TS U1137 ( .A(sumIn[65]), .B(n938), .Y(n1084) );
  OAI21XLTS U1138 ( .A0(n941), .A1(n947), .B0(n940), .Y(n939) );
  NAND2X1TS U1139 ( .A(n1088), .B(n942), .Y(n978) );
  NAND2X1TS U1140 ( .A(n1088), .B(n1084), .Y(n974) );
  AOI21X1TS U1141 ( .A0(n1088), .A1(n976), .B0(n942), .Y(n973) );
  XNOR2X1TS U1142 ( .A(sumIn[63]), .B(n943), .Y(n1113) );
  INVX2TS U1143 ( .A(n944), .Y(n965) );
  NOR3XLTS U1144 ( .A(n953), .B(n965), .C(n957), .Y(n949) );
  OAI21XLTS U1145 ( .A0(n949), .A1(n945), .B0(n948), .Y(n946) );
  OAI21XLTS U1146 ( .A0(n960), .A1(n950), .B0(n985), .Y(n951) );
  XNOR2X1TS U1147 ( .A(n952), .B(n951), .Y(n1094) );
  OAI21XLTS U1148 ( .A0(n965), .A1(n957), .B0(n962), .Y(n954) );
  OAI2BB2XLTS U1149 ( .B0(n1114), .B1(n968), .A0N(n1094), .A1N(n1097), .Y(n955) );
  OAI2BB1X1TS U1150 ( .A0N(n968), .A1N(n1114), .B0(n955), .Y(n972) );
  INVX2TS U1151 ( .A(n956), .Y(n1103) );
  NAND2X1TS U1152 ( .A(n1103), .B(n958), .Y(n959) );
  INVX2TS U1153 ( .A(n961), .Y(n1102) );
  NAND2X1TS U1154 ( .A(n962), .B(n1102), .Y(n964) );
  AOI222XLTS U1155 ( .A0(n967), .A1(n1106), .B0(n967), .B1(n966), .C0(n1106), 
        .C1(n965), .Y(n970) );
  NAND2X1TS U1156 ( .A(n1114), .B(n968), .Y(n969) );
  OAI211XLTS U1157 ( .A0(n1094), .A1(n1097), .B0(n970), .C0(n969), .Y(n971) );
  AOI22X1TS U1158 ( .A0(n974), .A1(n973), .B0(n972), .B1(n971), .Y(n975) );
  AOI21X1TS U1159 ( .A0(n1084), .A1(n976), .B0(n975), .Y(n977) );
  OAI211XLTS U1160 ( .A0(n1078), .A1(n1080), .B0(n978), .C0(n977), .Y(n979) );
  OAI2BB1X1TS U1161 ( .A0N(n1080), .A1N(n1078), .B0(n979), .Y(n980) );
  AOI222XLTS U1162 ( .A0(n981), .A1(n990), .B0(n981), .B1(n980), .C0(n990), 
        .C1(n980), .Y(n984) );
  NOR2XLTS U1163 ( .A(sumIn[77]), .B(n982), .Y(n987) );
  NOR2XLTS U1164 ( .A(n921), .B(n987), .Y(n983) );
  XNOR2X1TS U1165 ( .A(n983), .B(sumIn[78]), .Y(n1074) );
  AOI222XLTS U1166 ( .A0(n1073), .A1(n984), .B0(n1073), .B1(n1074), .C0(n984), 
        .C1(n1074), .Y(n988) );
  INVX2TS U1167 ( .A(n601), .Y(n1283) );
  INVX2TS U1168 ( .A(sumIn[82]), .Y(n991) );
  INVX2TS U1169 ( .A(n991), .Y(n1030) );
  INVX2TS U1170 ( .A(sumIn[81]), .Y(n992) );
  INVX2TS U1171 ( .A(n992), .Y(n1037) );
  INVX2TS U1172 ( .A(sumIn[80]), .Y(n1034) );
  INVX2TS U1173 ( .A(n1034), .Y(n1028) );
  NOR4XLTS U1174 ( .A(sumIn[83]), .B(n1030), .C(n1037), .D(n1028), .Y(n1009)
         );
  NOR2XLTS U1175 ( .A(sumIn[85]), .B(n1014), .Y(n1004) );
  INVX2TS U1176 ( .A(sumIn[89]), .Y(n1000) );
  INVX2TS U1177 ( .A(n1000), .Y(n1035) );
  NAND2X1TS U1178 ( .A(n1002), .B(n1035), .Y(n993) );
  INVX2TS U1179 ( .A(sumIn[93]), .Y(n994) );
  INVX2TS U1180 ( .A(n994), .Y(n1026) );
  INVX2TS U1181 ( .A(sumIn[92]), .Y(n995) );
  INVX2TS U1182 ( .A(n995), .Y(n1031) );
  INVX2TS U1183 ( .A(sumIn[91]), .Y(n1022) );
  INVX2TS U1184 ( .A(n1022), .Y(n1041) );
  INVX2TS U1185 ( .A(sumIn[90]), .Y(n1039) );
  INVX2TS U1186 ( .A(n1039), .Y(n1038) );
  NOR4XLTS U1187 ( .A(n1026), .B(n1031), .C(n1041), .D(n1038), .Y(n1018) );
  INVX2TS U1188 ( .A(sumIn[94]), .Y(n996) );
  INVX2TS U1189 ( .A(n996), .Y(n1017) );
  NOR2BX1TS U1190 ( .AN(n1018), .B(n1017), .Y(n1013) );
  INVX2TS U1191 ( .A(sumIn[95]), .Y(n997) );
  INVX2TS U1192 ( .A(n997), .Y(n1012) );
  NOR2BX1TS U1193 ( .AN(n1013), .B(n1012), .Y(n1007) );
  INVX2TS U1194 ( .A(sumIn[99]), .Y(n998) );
  INVX2TS U1195 ( .A(n998), .Y(n1040) );
  NAND2X1TS U1196 ( .A(n1061), .B(n1040), .Y(n999) );
  XNOR2X1TS U1197 ( .A(sumIn[97]), .B(n999), .Y(n1060) );
  INVX2TS U1198 ( .A(n1000), .Y(n1065) );
  NOR2XLTS U1199 ( .A(sumIn[87]), .B(n1002), .Y(n1066) );
  OAI21XLTS U1200 ( .A0(n1066), .A1(n1001), .B0(sumIn[88]), .Y(n1003) );
  OAI21XLTS U1201 ( .A0(sumIn[88]), .A1(n1001), .B0(n1003), .Y(n1077) );
  NOR2XLTS U1202 ( .A(n1000), .B(n1004), .Y(n1005) );
  CLKBUFX2TS U1203 ( .A(n1040), .Y(n1010) );
  INVX2TS U1204 ( .A(n1010), .Y(n1025) );
  INVX2TS U1205 ( .A(n1010), .Y(n1023) );
  OAI21XLTS U1206 ( .A0(n1007), .A1(n1023), .B0(sumIn[96]), .Y(n1006) );
  OAI31XLTS U1207 ( .A0(n1007), .A1(sumIn[96]), .A2(n1025), .B0(n1006), .Y(
        n1081) );
  OAI21XLTS U1208 ( .A0(n1009), .A1(n1001), .B0(sumIn[84]), .Y(n1008) );
  OAI31XLTS U1209 ( .A0(n1009), .A1(sumIn[84]), .A2(n1001), .B0(n1008), .Y(
        n1086) );
  OAI21XLTS U1210 ( .A0(n1013), .A1(n1025), .B0(n1012), .Y(n1011) );
  NAND2X1TS U1211 ( .A(n1014), .B(n1035), .Y(n1015) );
  XNOR2X1TS U1212 ( .A(sumIn[85]), .B(n1015), .Y(n1054) );
  OAI21XLTS U1213 ( .A0(n1018), .A1(n1025), .B0(n1017), .Y(n1016) );
  AOI21X1TS U1214 ( .A0(n1019), .A1(n1083), .B0(n1087), .Y(n1020) );
  NAND2X1TS U1215 ( .A(n1086), .B(n1020), .Y(n1056) );
  NAND2X1TS U1216 ( .A(n1086), .B(n1054), .Y(n1051) );
  AOI21X1TS U1217 ( .A0(n1086), .A1(n1053), .B0(n1020), .Y(n1050) );
  INVX2TS U1218 ( .A(n1022), .Y(n1043) );
  NOR3XLTS U1219 ( .A(n1031), .B(n1043), .C(n1038), .Y(n1027) );
  OAI21XLTS U1220 ( .A0(n1027), .A1(n1023), .B0(n1026), .Y(n1024) );
  OAI21XLTS U1221 ( .A0(n1037), .A1(n1028), .B0(n1065), .Y(n1029) );
  XNOR2X1TS U1222 ( .A(n1030), .B(n1029), .Y(n1099) );
  OAI21XLTS U1223 ( .A0(n1043), .A1(n1038), .B0(n1040), .Y(n1032) );
  OAI2BB2XLTS U1224 ( .B0(n1090), .B1(n1092), .A0N(n1099), .A1N(n1098), .Y(
        n1033) );
  OAI2BB1X1TS U1225 ( .A0N(n1092), .A1N(n1090), .B0(n1033), .Y(n1049) );
  INVX2TS U1226 ( .A(n1034), .Y(n1110) );
  NAND2X1TS U1227 ( .A(n1035), .B(n1110), .Y(n1036) );
  XNOR2X1TS U1228 ( .A(n1037), .B(n1036), .Y(n1104) );
  INVX2TS U1229 ( .A(n1039), .Y(n1109) );
  NAND2X1TS U1230 ( .A(n1040), .B(n1109), .Y(n1042) );
  XNOR2X1TS U1231 ( .A(n1042), .B(n1041), .Y(n1105) );
  AOI222XLTS U1232 ( .A0(n1045), .A1(n1044), .B0(n1045), .B1(n1043), .C0(n1044), .C1(n1105), .Y(n1047) );
  NAND2X1TS U1233 ( .A(n1090), .B(n1092), .Y(n1046) );
  OAI211XLTS U1234 ( .A0(n1099), .A1(n1098), .B0(n1047), .C0(n1046), .Y(n1048)
         );
  AOI22X1TS U1235 ( .A0(n1051), .A1(n1050), .B0(n1049), .B1(n1048), .Y(n1052)
         );
  AOI21X1TS U1236 ( .A0(n1054), .A1(n1053), .B0(n1052), .Y(n1055) );
  OAI211XLTS U1237 ( .A0(n1081), .A1(n1058), .B0(n1056), .C0(n1055), .Y(n1057)
         );
  OAI2BB1X1TS U1238 ( .A0N(n1058), .A1N(n1081), .B0(n1057), .Y(n1059) );
  AOI222XLTS U1239 ( .A0(n1060), .A1(n1070), .B0(n1060), .B1(n1059), .C0(n1070), .C1(n1059), .Y(n1064) );
  NOR2XLTS U1240 ( .A(sumIn[97]), .B(n1061), .Y(n1067) );
  NOR2XLTS U1241 ( .A(n998), .B(n1067), .Y(n1062) );
  AOI222XLTS U1242 ( .A0(n1077), .A1(n1064), .B0(n1077), .B1(n1063), .C0(n1064), .C1(n1063), .Y(n1068) );
  INVX2TS U1243 ( .A(n602), .Y(n1284) );
  NOR2BX1TS U1244 ( .AN(n1072), .B(n1071), .Y(n1191) );
  INVX2TS U1245 ( .A(n602), .Y(n1091) );
  INVX2TS U1246 ( .A(n601), .Y(n1095) );
  NAND2X1TS U1247 ( .A(n1142), .B(n1140), .Y(n1118) );
  OAI21XLTS U1248 ( .A0(n1157), .A1(n1159), .B0(n1152), .Y(n1111) );
  OAI2BB2XLTS U1249 ( .B0(n1153), .B1(n1111), .A0N(n1157), .A1N(n1159), .Y(
        n1112) );
  AOI222XLTS U1250 ( .A0(n1151), .A1(n1149), .B0(n1151), .B1(n1112), .C0(n1149), .C1(n1112), .Y(n1115) );
  AOI222XLTS U1251 ( .A0(n1168), .A1(n1115), .B0(n1168), .B1(n1170), .C0(n1115), .C1(n1170), .Y(n1116) );
  OAI211XLTS U1252 ( .A0(n1172), .A1(n1119), .B0(n1118), .C0(n1117), .Y(n1120)
         );
  OAI21XLTS U1253 ( .A0(n1142), .A1(n1140), .B0(n1120), .Y(n1121) );
  AOI222XLTS U1254 ( .A0(n1135), .A1(n1136), .B0(n1135), .B1(n1121), .C0(n1136), .C1(n1121), .Y(n1122) );
  AOI222XLTS U1255 ( .A0(n1129), .A1(n1123), .B0(n1129), .B1(n1122), .C0(n1123), .C1(n1122), .Y(n1124) );
  OAI21XLTS U1256 ( .A0(n1131), .A1(n1132), .B0(n1124), .Y(n1128) );
  NAND2X1TS U1257 ( .A(n1131), .B(n1132), .Y(n1127) );
  AOI31XLTS U1258 ( .A0(n1191), .A1(n1128), .A2(n1127), .B0(n1192), .Y(n1282)
         );
  INVX2TS U1259 ( .A(n1282), .Y(n1141) );
  NOR2BX1TS U1260 ( .AN(n1132), .B(n1131), .Y(n1265) );
  INVX2TS U1261 ( .A(n1144), .Y(n1180) );
  INVX2TS U1262 ( .A(n1144), .Y(n1286) );
  INVX2TS U1263 ( .A(n1282), .Y(n1292) );
  INVX2TS U1264 ( .A(n1282), .Y(n1285) );
  OAI21XLTS U1265 ( .A0(n1222), .A1(n1223), .B0(n1219), .Y(n1162) );
  OAI2BB2XLTS U1266 ( .B0(n1221), .B1(n1162), .A0N(n1222), .A1N(n1223), .Y(
        n1167) );
  AOI222XLTS U1267 ( .A0(n1213), .A1(n1167), .B0(n1213), .B1(n1215), .C0(n1167), .C1(n1215), .Y(n1171) );
  AOI222XLTS U1268 ( .A0(n1210), .A1(n1171), .B0(n1210), .B1(n1208), .C0(n1171), .C1(n1208), .Y(n1177) );
  NOR2XLTS U1269 ( .A(n1202), .B(n1204), .Y(n1174) );
  NOR2XLTS U1270 ( .A(n1206), .B(n1174), .Y(n1176) );
  AOI21X1TS U1271 ( .A0(n1204), .A1(n1202), .B0(n1179), .Y(n1187) );
  NAND2X1TS U1272 ( .A(n1189), .B(n1198), .Y(n1183) );
  NAND2X1TS U1273 ( .A(n1200), .B(n1183), .Y(n1184) );
  OAI2BB1X1TS U1274 ( .A0N(n1201), .A1N(n1187), .B0(n1186), .Y(n1188) );
  OAI21XLTS U1275 ( .A0(n1198), .A1(n1189), .B0(n1188), .Y(n1190) );
  AOI222XLTS U1276 ( .A0(n1265), .A1(n1268), .B0(n1265), .B1(n1190), .C0(n1268), .C1(n1190), .Y(n1193) );
  AOI21X1TS U1277 ( .A0(n1194), .A1(n1193), .B0(n1279), .Y(n1195) );
  INVX2TS U1278 ( .A(n1195), .Y(n1199) );
  INVX2TS U1279 ( .A(n1199), .Y(n1294) );
  INVX2TS U1280 ( .A(n1195), .Y(n1266) );
  INVX2TS U1281 ( .A(n1246), .Y(n1232) );
  OAI21XLTS U1282 ( .A0(n1219), .A1(n1266), .B0(n1218), .Y(n1220) );
  CLKBUFX2TS U1283 ( .A(n1225), .Y(n1246) );
  AOI222XLTS U1284 ( .A0(n1230), .A1(n1229), .B0(n1230), .B1(n1228), .C0(n1229), .C1(n1228), .Y(n1238) );
  OA21XLTS U1285 ( .A0(n1238), .A1(n1239), .B0(n1235), .Y(n1237) );
  NOR2XLTS U1286 ( .A(n1242), .B(n1241), .Y(n1236) );
  AOI211XLTS U1287 ( .A0(n1239), .A1(n1238), .B0(n1237), .C0(n1236), .Y(n1240)
         );
  AOI21X1TS U1288 ( .A0(n1242), .A1(n1241), .B0(n1240), .Y(n1251) );
  AOI21X1TS U1289 ( .A0(n1244), .A1(n1246), .B0(n1249), .Y(n1245) );
  OAI21XLTS U1290 ( .A0(n1247), .A1(n1246), .B0(n1245), .Y(n1248) );
  OAI2BB1X1TS U1291 ( .A0N(n1252), .A1N(n1251), .B0(n1250), .Y(n1253) );
  OAI21XLTS U1292 ( .A0(n1255), .A1(n1254), .B0(n1253), .Y(n1259) );
  AOI222XLTS U1293 ( .A0(n1260), .A1(n1259), .B0(n1260), .B1(n1258), .C0(n1259), .C1(n1258), .Y(n1261) );
  OAI2BB1X1TS U1294 ( .A0N(n1264), .A1N(n1263), .B0(n1261), .Y(n1262) );
  NOR2BX1TS U1295 ( .AN(n1270), .B(n1269), .Y(n1272) );
  NAND2X1TS U1296 ( .A(n1274), .B(n1273), .Y(n1271) );
  OAI2BB2XLTS U1297 ( .B0(n1274), .B1(n1273), .A0N(n1272), .A1N(n1271), .Y(
        n1280) );
  OAI31X1TS U1298 ( .A0(n1281), .A1(n1280), .A2(n1279), .B0(n1278), .Y(
        result[3]) );
  AOI22X1TS U1299 ( .A0(n1285), .A1(n1284), .B0(n1283), .B1(n1282), .Y(n1291)
         );
  NOR2XLTS U1300 ( .A(result[3]), .B(n1199), .Y(result[2]) );
  AOI22X1TS U1301 ( .A0(n1293), .A1(n1288), .B0(n1287), .B1(n1286), .Y(n1289)
         );
  AOI22X1TS U1302 ( .A0(n1232), .A1(result[3]), .B0(result[2]), .B1(n1289), 
        .Y(n1290) );
  OAI31X1TS U1303 ( .A0(n1294), .A1(result[3]), .A2(n1291), .B0(n1290), .Y(
        result[0]) );
  AOI221XLTS U1304 ( .A0(n1294), .A1(n1293), .B0(n1196), .B1(n1292), .C0(
        result[3]), .Y(result[1]) );
endmodule

